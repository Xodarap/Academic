library verilog;
use verilog.vl_types.all;
entity tb_shifter1 is
end tb_shifter1;
