library verilog;
use verilog.vl_types.all;
entity mem_system_hier_tb is
end mem_system_hier_tb;
