library verilog;
use verilog.vl_types.all;
entity tb_shifter is
end tb_shifter;
