library verilog;
use verilog.vl_types.all;
entity tb_cond_set is
end tb_cond_set;
