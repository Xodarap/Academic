library verilog;
use verilog.vl_types.all;
entity tb_rf_hier is
end tb_rf_hier;
