library verilog;
use verilog.vl_types.all;
entity rf_bypass_bench is
end rf_bypass_bench;
