library verilog;
use verilog.vl_types.all;
entity tb_fetch is
end tb_fetch;
