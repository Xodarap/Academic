library verilog;
use verilog.vl_types.all;
entity tb_control is
end tb_control;
