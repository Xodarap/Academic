library verilog;
use verilog.vl_types.all;
entity proc_hier is
end proc_hier;
