library verilog;
use verilog.vl_types.all;
entity seq_detect_bench is
end seq_detect_bench;
