library verilog;
use verilog.vl_types.all;
entity tb_onebitreg is
end tb_onebitreg;
