library verilog;
use verilog.vl_types.all;
entity mem_system_randbench is
end mem_system_randbench;
