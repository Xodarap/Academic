
module xor2_7 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_6 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module nand2_11 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_10 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_9 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module xor2_5 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_4 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module nand2_8 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_7 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_6 ( in1, in2, out );
  input in1, in2;
  output out;


  NAND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_3 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_2 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module nand2_5 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_4 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_3 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module xor2_1 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module xor2_0 ( in1, in2, out );
  input in1, in2;
  output out;


  XOR2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module nand2_2 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_1 ( in1, in2, out );
  input in1, in2;
  output out;
  wire   n1;

  AND2X1 U1 ( .A(in2), .B(in1), .Y(n1) );
  INVX1 U2 ( .A(n1), .Y(out) );
endmodule


module nand2_0 ( in1, in2, out );
  input in1, in2;
  output out;


  NAND2X1 U1 ( .A(in2), .B(in1), .Y(out) );
endmodule


module dff_0 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_1 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_2 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_3 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  OR2X1 U3 ( .A(n3), .B(rst), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
  INVX1 U5 ( .A(d), .Y(n3) );
endmodule


module fulladder1_3 ( A, B, Cin, S, Cout );
  input A, B, Cin;
  output S, Cout;
  wire   x1_out, n1_out, n2_out;

  xor2_7 x1 ( .in1(A), .in2(B), .out(x1_out) );
  xor2_6 x2 ( .in1(x1_out), .in2(Cin), .out(S) );
  nand2_11 n1 ( .in1(A), .in2(B), .out(n1_out) );
  nand2_10 n2 ( .in1(x1_out), .in2(Cin), .out(n2_out) );
  nand2_9 n3 ( .in1(n2_out), .in2(n1_out), .out(Cout) );
endmodule


module fulladder1_2 ( A, B, Cin, S, Cout );
  input A, B, Cin;
  output S, Cout;
  wire   x1_out, n1_out, n2_out;

  xor2_5 x1 ( .in1(A), .in2(B), .out(x1_out) );
  xor2_4 x2 ( .in1(x1_out), .in2(Cin), .out(S) );
  nand2_8 n1 ( .in1(A), .in2(B), .out(n1_out) );
  nand2_7 n2 ( .in1(x1_out), .in2(Cin), .out(n2_out) );
  nand2_6 n3 ( .in1(n2_out), .in2(n1_out), .out(Cout) );
endmodule


module fulladder1_1 ( A, B, Cin, S, Cout );
  input A, B, Cin;
  output S, Cout;
  wire   x1_out, n1_out, n2_out;

  xor2_3 x1 ( .in1(A), .in2(B), .out(x1_out) );
  xor2_2 x2 ( .in1(x1_out), .in2(Cin), .out(S) );
  nand2_5 n1 ( .in1(A), .in2(B), .out(n1_out) );
  nand2_4 n2 ( .in1(x1_out), .in2(Cin), .out(n2_out) );
  nand2_3 n3 ( .in1(n2_out), .in2(n1_out), .out(Cout) );
endmodule


module fulladder1_0 ( A, B, Cin, S, Cout );
  input A, B, Cin;
  output S, Cout;
  wire   x1_out, n1_out, n2_out;

  xor2_1 x1 ( .in1(A), .in2(B), .out(x1_out) );
  xor2_0 x2 ( .in1(x1_out), .in2(Cin), .out(S) );
  nand2_2 n1 ( .in1(A), .in2(B), .out(n1_out) );
  nand2_1 n2 ( .in1(x1_out), .in2(Cin), .out(n2_out) );
  nand2_0 n3 ( .in1(n2_out), .in2(n1_out), .out(Cout) );
endmodule


module onebitreg_0 ( readdata, clk, rst, writedata, write );
  input clk, rst, writedata, write;
  output readdata;
  wire   n3, n1, n2, n4;

  AOI22X1 U3 ( .A(readdata), .B(n4), .C(writedata), .D(write), .Y(n3) );
  dff_0 data ( .q(readdata), .d(n2), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(write), .Y(n4) );
  BUFX2 U2 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
endmodule


module onebitreg_1 ( readdata, clk, rst, writedata, write );
  input clk, rst, writedata, write;
  output readdata;
  wire   n1, n2, n4, n5;

  AOI22X1 U3 ( .A(readdata), .B(n4), .C(writedata), .D(write), .Y(n5) );
  dff_1 data ( .q(readdata), .d(n2), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(write), .Y(n4) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
endmodule


module onebitreg_2 ( readdata, clk, rst, writedata, write );
  input clk, rst, writedata, write;
  output readdata;
  wire   n1, n2, n4, n5;

  AOI22X1 U3 ( .A(readdata), .B(n4), .C(writedata), .D(write), .Y(n5) );
  dff_2 data ( .q(readdata), .d(n2), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(write), .Y(n4) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
endmodule


module onebitreg_3 ( readdata, clk, rst, writedata, write );
  input clk, rst, writedata, write;
  output readdata;
  wire   n1, n2, n4, n5;

  AOI22X1 U3 ( .A(readdata), .B(n4), .C(writedata), .D(write), .Y(n5) );
  dff_3 data ( .q(readdata), .d(n2), .clk(clk), .rst(rst) );
  INVX1 U1 ( .A(write), .Y(n4) );
  BUFX2 U2 ( .A(n5), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n2) );
endmodule


module dff_200 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_201 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_202 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_203 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_204 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_205 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_206 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_207 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_208 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_209 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_210 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_211 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_212 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_213 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_214 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_215 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_216 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_217 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_218 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_219 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_220 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_221 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_222 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_223 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_224 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_225 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_226 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_227 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_228 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_229 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_230 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_231 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_232 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_233 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_234 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_235 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_236 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_237 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_238 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_239 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_240 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_241 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_242 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_243 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_244 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_245 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_246 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_247 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_248 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_249 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_250 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_251 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_252 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_253 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_254 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_255 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_256 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_257 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_258 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_259 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_260 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_261 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_262 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_263 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_136 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_137 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_138 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_139 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_140 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_141 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_142 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_143 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_144 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_145 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_146 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_147 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_148 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_149 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_150 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_151 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_152 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_153 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_154 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_155 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_156 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_157 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_158 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_159 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_160 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_161 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_162 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_163 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_164 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_165 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_166 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_167 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_168 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_169 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_170 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_171 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_172 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_173 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_174 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_175 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_176 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_177 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_178 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_179 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_180 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_181 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_182 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_183 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_184 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_185 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_186 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_187 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_188 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_189 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_190 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_191 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_192 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_193 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_194 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_195 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_196 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_197 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_198 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_199 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_72 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_73 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_74 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_75 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_76 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_77 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_78 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_79 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_80 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_81 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_82 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_83 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_84 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_85 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_86 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_87 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_88 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_89 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_90 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_91 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_92 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_93 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_94 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_95 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_96 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_97 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_98 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_99 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_100 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_101 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_102 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_103 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_104 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_105 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_106 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_107 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_108 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_109 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_110 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_111 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_112 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_113 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_114 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_115 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_116 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_117 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_118 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_119 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_120 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_121 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_122 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_123 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_124 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_125 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_126 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_127 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_128 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_129 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_130 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_131 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_132 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_133 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_134 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_135 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_8 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_9 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_10 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_11 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_12 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_13 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_14 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_15 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_16 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_17 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_18 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_19 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_20 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_21 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_22 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_23 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_24 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_25 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_26 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_27 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_28 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_29 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_30 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_31 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_32 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_33 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_34 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_35 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_36 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_37 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_38 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_39 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_40 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_41 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_42 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_43 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_44 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_45 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_46 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_47 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_48 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_49 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_50 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_51 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_52 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_53 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_54 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_55 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_56 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_57 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_58 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_59 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_60 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_61 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_62 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_63 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_64 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_65 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_66 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_67 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_68 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_69 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_70 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_71 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module fulladder2_1 ( .A({\A<1> , \A<0> }), .B({\B<1> , \B<0> }), .SUM({
        \SUM<1> , \SUM<0> }) );
  input \A<1> , \A<0> , \B<1> , \B<0> ;
  output \SUM<1> , \SUM<0> ;
  wire   c1;

  fulladder1_3 add0 ( .A(\A<0> ), .B(\B<0> ), .Cin(1'b0), .S(\SUM<0> ), .Cout(
        c1) );
  fulladder1_2 add1 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .S(\SUM<1> ), .Cout()
         );
endmodule


module fulladder2_0 ( .A({\A<1> , \A<0> }), .B({\B<1> , \B<0> }), .SUM({
        \SUM<1> , \SUM<0> }) );
  input \A<1> , \A<0> , \B<1> , \B<0> ;
  output \SUM<1> , \SUM<0> ;
  wire   c1;

  fulladder1_1 add0 ( .A(\A<0> ), .B(\B<0> ), .Cin(1'b0), .S(\SUM<0> ), .Cout(
        c1) );
  fulladder1_0 add1 ( .A(\A<1> ), .B(\B<1> ), .Cin(c1), .S(\SUM<1> ), .Cout()
         );
endmodule


module counter5 ( push, pop, rst, clk, .currentState({\currentState<3> , 
        \currentState<2> , \currentState<1> , \currentState<0> }) );
  input push, pop, rst, clk;
  output \currentState<3> , \currentState<2> , \currentState<1> ,
         \currentState<0> ;
  wire   \nextReg<2> , n17, n21, n22, n23, n24, n26, n27, n28, n29, n30, n31,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n25, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  FAX1 U11 ( .A(n34), .B(\currentState<3> ), .C(n3), .YC(), .YS(n17) );
  OAI21X1 U14 ( .A(n2), .B(n22), .C(n23), .Y(\nextReg<2> ) );
  FAX1 U15 ( .A(\currentState<2> ), .B(n34), .C(n21), .YC(), .YS(n22) );
  OAI21X1 U16 ( .A(n34), .B(n1), .C(n26), .Y(n21) );
  OAI21X1 U17 ( .A(n4), .B(n38), .C(\currentState<1> ), .Y(n26) );
  FAX1 U19 ( .A(\currentState<1> ), .B(n38), .C(n1), .YC(), .YS(n27) );
  XNOR2X1 U22 ( .A(\currentState<0> ), .B(n28), .Y(n29) );
  OAI21X1 U23 ( .A(pop), .B(n39), .C(n34), .Y(n28) );
  NAND3X1 U25 ( .A(n31), .B(n34), .C(\currentState<2> ), .Y(n24) );
  NAND3X1 U26 ( .A(n31), .B(n40), .C(n38), .Y(n30) );
  NOR3X1 U28 ( .A(\currentState<1> ), .B(\currentState<3> ), .C(
        \currentState<0> ), .Y(n31) );
  onebitreg_0 \state[0]  ( .readdata(\currentState<0> ), .clk(clk), .rst(n35), 
        .writedata(n16), .write(1'b1) );
  onebitreg_1 \state[1]  ( .readdata(\currentState<1> ), .clk(clk), .rst(n35), 
        .writedata(n19), .write(1'b1) );
  onebitreg_2 \state[2]  ( .readdata(\currentState<2> ), .clk(clk), .rst(n35), 
        .writedata(\nextReg<2> ), .write(1'b1) );
  onebitreg_3 \state[3]  ( .readdata(\currentState<3> ), .clk(clk), .rst(n35), 
        .writedata(n6), .write(1'b1) );
  AND2X2 U3 ( .A(n10), .B(n14), .Y(n3) );
  AND2X2 U4 ( .A(\currentState<0> ), .B(n28), .Y(n4) );
  INVX2 U5 ( .A(n4), .Y(n1) );
  INVX2 U6 ( .A(n36), .Y(n35) );
  OR2X1 U7 ( .A(n20), .B(n35), .Y(n23) );
  OR2X1 U8 ( .A(n2), .B(n17), .Y(n5) );
  OR2X1 U9 ( .A(n32), .B(n12), .Y(n2) );
  INVX4 U10 ( .A(n33), .Y(n34) );
  AND2X2 U12 ( .A(pop), .B(n39), .Y(n33) );
  AND2X2 U13 ( .A(n37), .B(n34), .Y(n13) );
  INVX1 U18 ( .A(push), .Y(n39) );
  INVX1 U20 ( .A(n5), .Y(n6) );
  AND2X2 U21 ( .A(n38), .B(n21), .Y(n7) );
  INVX1 U24 ( .A(n7), .Y(n8) );
  AND2X2 U27 ( .A(n40), .B(n8), .Y(n9) );
  INVX1 U29 ( .A(n9), .Y(n10) );
  BUFX2 U30 ( .A(n30), .Y(n11) );
  INVX1 U31 ( .A(n34), .Y(n38) );
  OR2X1 U32 ( .A(n25), .B(rst), .Y(n12) );
  INVX1 U33 ( .A(n13), .Y(n14) );
  OR2X1 U34 ( .A(n2), .B(n29), .Y(n15) );
  INVX1 U35 ( .A(n15), .Y(n16) );
  OR2X1 U36 ( .A(n27), .B(n2), .Y(n18) );
  INVX1 U37 ( .A(n18), .Y(n19) );
  BUFX2 U38 ( .A(n24), .Y(n20) );
  INVX1 U39 ( .A(\currentState<2> ), .Y(n40) );
  INVX1 U40 ( .A(n21), .Y(n37) );
  INVX1 U41 ( .A(n20), .Y(n25) );
  INVX1 U42 ( .A(n11), .Y(n32) );
  INVX1 U43 ( .A(rst), .Y(n36) );
endmodule


module dff_6 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_7 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_4 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module dff_5 ( q, d, clk, rst );
  input d, clk, rst;
  output q;
  wire   n1, n2, n3;

  DFFPOSX1 state_reg ( .D(n2), .CLK(clk), .Q(q) );
  INVX1 U3 ( .A(d), .Y(n3) );
  OR2X1 U4 ( .A(rst), .B(n3), .Y(n1) );
  INVX1 U5 ( .A(n1), .Y(n2) );
endmodule


module fifo ( .data_out({\data_out<63> , \data_out<62> , \data_out<61> , 
        \data_out<60> , \data_out<59> , \data_out<58> , \data_out<57> , 
        \data_out<56> , \data_out<55> , \data_out<54> , \data_out<53> , 
        \data_out<52> , \data_out<51> , \data_out<50> , \data_out<49> , 
        \data_out<48> , \data_out<47> , \data_out<46> , \data_out<45> , 
        \data_out<44> , \data_out<43> , \data_out<42> , \data_out<41> , 
        \data_out<40> , \data_out<39> , \data_out<38> , \data_out<37> , 
        \data_out<36> , \data_out<35> , \data_out<34> , \data_out<33> , 
        \data_out<32> , \data_out<31> , \data_out<30> , \data_out<29> , 
        \data_out<28> , \data_out<27> , \data_out<26> , \data_out<25> , 
        \data_out<24> , \data_out<23> , \data_out<22> , \data_out<21> , 
        \data_out<20> , \data_out<19> , \data_out<18> , \data_out<17> , 
        \data_out<16> , \data_out<15> , \data_out<14> , \data_out<13> , 
        \data_out<12> , \data_out<11> , \data_out<10> , \data_out<9> , 
        \data_out<8> , \data_out<7> , \data_out<6> , \data_out<5> , 
        \data_out<4> , \data_out<3> , \data_out<2> , \data_out<1> , 
        \data_out<0> }), fifo_empty, fifo_full, data_out_valid, err, 
    .data_in({\data_in<63> , \data_in<62> , \data_in<61> , \data_in<60> , 
        \data_in<59> , \data_in<58> , \data_in<57> , \data_in<56> , 
        \data_in<55> , \data_in<54> , \data_in<53> , \data_in<52> , 
        \data_in<51> , \data_in<50> , \data_in<49> , \data_in<48> , 
        \data_in<47> , \data_in<46> , \data_in<45> , \data_in<44> , 
        \data_in<43> , \data_in<42> , \data_in<41> , \data_in<40> , 
        \data_in<39> , \data_in<38> , \data_in<37> , \data_in<36> , 
        \data_in<35> , \data_in<34> , \data_in<33> , \data_in<32> , 
        \data_in<31> , \data_in<30> , \data_in<29> , \data_in<28> , 
        \data_in<27> , \data_in<26> , \data_in<25> , \data_in<24> , 
        \data_in<23> , \data_in<22> , \data_in<21> , \data_in<20> , 
        \data_in<19> , \data_in<18> , \data_in<17> , \data_in<16> , 
        \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> , 
        \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> , \data_in<7> , 
        \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> , \data_in<2> , 
        \data_in<1> , \data_in<0> }), data_in_valid, pop_fifo, clk, rst );
  input \data_in<63> , \data_in<62> , \data_in<61> , \data_in<60> ,
         \data_in<59> , \data_in<58> , \data_in<57> , \data_in<56> ,
         \data_in<55> , \data_in<54> , \data_in<53> , \data_in<52> ,
         \data_in<51> , \data_in<50> , \data_in<49> , \data_in<48> ,
         \data_in<47> , \data_in<46> , \data_in<45> , \data_in<44> ,
         \data_in<43> , \data_in<42> , \data_in<41> , \data_in<40> ,
         \data_in<39> , \data_in<38> , \data_in<37> , \data_in<36> ,
         \data_in<35> , \data_in<34> , \data_in<33> , \data_in<32> ,
         \data_in<31> , \data_in<30> , \data_in<29> , \data_in<28> ,
         \data_in<27> , \data_in<26> , \data_in<25> , \data_in<24> ,
         \data_in<23> , \data_in<22> , \data_in<21> , \data_in<20> ,
         \data_in<19> , \data_in<18> , \data_in<17> , \data_in<16> ,
         \data_in<15> , \data_in<14> , \data_in<13> , \data_in<12> ,
         \data_in<11> , \data_in<10> , \data_in<9> , \data_in<8> ,
         \data_in<7> , \data_in<6> , \data_in<5> , \data_in<4> , \data_in<3> ,
         \data_in<2> , \data_in<1> , \data_in<0> , data_in_valid, pop_fifo,
         clk, rst;
  output \data_out<63> , \data_out<62> , \data_out<61> , \data_out<60> ,
         \data_out<59> , \data_out<58> , \data_out<57> , \data_out<56> ,
         \data_out<55> , \data_out<54> , \data_out<53> , \data_out<52> ,
         \data_out<51> , \data_out<50> , \data_out<49> , \data_out<48> ,
         \data_out<47> , \data_out<46> , \data_out<45> , \data_out<44> ,
         \data_out<43> , \data_out<42> , \data_out<41> , \data_out<40> ,
         \data_out<39> , \data_out<38> , \data_out<37> , \data_out<36> ,
         \data_out<35> , \data_out<34> , \data_out<33> , \data_out<32> ,
         \data_out<31> , \data_out<30> , \data_out<29> , \data_out<28> ,
         \data_out<27> , \data_out<26> , \data_out<25> , \data_out<24> ,
         \data_out<23> , \data_out<22> , \data_out<21> , \data_out<20> ,
         \data_out<19> , \data_out<18> , \data_out<17> , \data_out<16> ,
         \data_out<15> , \data_out<14> , \data_out<13> , \data_out<12> ,
         \data_out<11> , \data_out<10> , \data_out<9> , \data_out<8> ,
         \data_out<7> , \data_out<6> , \data_out<5> , \data_out<4> ,
         \data_out<3> , \data_out<2> , \data_out<1> , \data_out<0> ,
         fifo_empty, fifo_full, data_out_valid, err;
  wire   \fifo0<63> , \fifo0<62> , \fifo0<61> , \fifo0<60> , \fifo0<59> ,
         \fifo0<58> , \fifo0<57> , \fifo0<56> , \fifo0<55> , \fifo0<54> ,
         \fifo0<53> , \fifo0<52> , \fifo0<51> , \fifo0<50> , \fifo0<49> ,
         \fifo0<48> , \fifo0<47> , \fifo0<46> , \fifo0<45> , \fifo0<44> ,
         \fifo0<43> , \fifo0<42> , \fifo0<41> , \fifo0<40> , \fifo0<39> ,
         \fifo0<38> , \fifo0<37> , \fifo0<36> , \fifo0<35> , \fifo0<34> ,
         \fifo0<33> , \fifo0<32> , \fifo0<31> , \fifo0<30> , \fifo0<29> ,
         \fifo0<28> , \fifo0<27> , \fifo0<26> , \fifo0<25> , \fifo0<24> ,
         \fifo0<23> , \fifo0<22> , \fifo0<21> , \fifo0<20> , \fifo0<19> ,
         \fifo0<18> , \fifo0<17> , \fifo0<16> , \fifo0<15> , \fifo0<14> ,
         \fifo0<13> , \fifo0<12> , \fifo0<11> , \fifo0<10> , \fifo0<9> ,
         \fifo0<8> , \fifo0<7> , \fifo0<6> , \fifo0<5> , \fifo0<4> ,
         \fifo0<3> , \fifo0<2> , \fifo0<1> , \fifo0<0> , \fifo_next0<63> ,
         \fifo_next0<62> , \fifo_next0<61> , \fifo_next0<60> ,
         \fifo_next0<59> , \fifo_next0<58> , \fifo_next0<57> ,
         \fifo_next0<56> , \fifo_next0<55> , \fifo_next0<54> ,
         \fifo_next0<53> , \fifo_next0<52> , \fifo_next0<51> ,
         \fifo_next0<50> , \fifo_next0<49> , \fifo_next0<48> ,
         \fifo_next0<47> , \fifo_next0<46> , \fifo_next0<45> ,
         \fifo_next0<44> , \fifo_next0<43> , \fifo_next0<42> ,
         \fifo_next0<41> , \fifo_next0<40> , \fifo_next0<39> ,
         \fifo_next0<38> , \fifo_next0<37> , \fifo_next0<36> ,
         \fifo_next0<35> , \fifo_next0<34> , \fifo_next0<33> ,
         \fifo_next0<32> , \fifo_next0<31> , \fifo_next0<30> ,
         \fifo_next0<29> , \fifo_next0<28> , \fifo_next0<27> ,
         \fifo_next0<26> , \fifo_next0<25> , \fifo_next0<24> ,
         \fifo_next0<23> , \fifo_next0<22> , \fifo_next0<21> ,
         \fifo_next0<20> , \fifo_next0<19> , \fifo_next0<18> ,
         \fifo_next0<17> , \fifo_next0<16> , \fifo_next0<15> ,
         \fifo_next0<14> , \fifo_next0<13> , \fifo_next0<12> ,
         \fifo_next0<11> , \fifo_next0<10> , \fifo_next0<9> , \fifo_next0<8> ,
         \fifo_next0<7> , \fifo_next0<6> , \fifo_next0<5> , \fifo_next0<4> ,
         \fifo_next0<3> , \fifo_next0<2> , \fifo_next0<1> , \fifo_next0<0> ,
         \fifo1<63> , \fifo1<62> , \fifo1<61> , \fifo1<60> , \fifo1<59> ,
         \fifo1<58> , \fifo1<57> , \fifo1<56> , \fifo1<55> , \fifo1<54> ,
         \fifo1<53> , \fifo1<52> , \fifo1<51> , \fifo1<50> , \fifo1<49> ,
         \fifo1<48> , \fifo1<47> , \fifo1<46> , \fifo1<45> , \fifo1<44> ,
         \fifo1<43> , \fifo1<42> , \fifo1<41> , \fifo1<40> , \fifo1<39> ,
         \fifo1<38> , \fifo1<37> , \fifo1<36> , \fifo1<35> , \fifo1<34> ,
         \fifo1<33> , \fifo1<32> , \fifo1<31> , \fifo1<30> , \fifo1<29> ,
         \fifo1<28> , \fifo1<27> , \fifo1<26> , \fifo1<25> , \fifo1<24> ,
         \fifo1<23> , \fifo1<22> , \fifo1<21> , \fifo1<20> , \fifo1<19> ,
         \fifo1<18> , \fifo1<17> , \fifo1<16> , \fifo1<15> , \fifo1<14> ,
         \fifo1<13> , \fifo1<12> , \fifo1<11> , \fifo1<10> , \fifo1<9> ,
         \fifo1<8> , \fifo1<7> , \fifo1<6> , \fifo1<5> , \fifo1<4> ,
         \fifo1<3> , \fifo1<2> , \fifo1<1> , \fifo1<0> , \fifo_next1<63> ,
         \fifo_next1<62> , \fifo_next1<61> , \fifo_next1<60> ,
         \fifo_next1<59> , \fifo_next1<58> , \fifo_next1<57> ,
         \fifo_next1<56> , \fifo_next1<55> , \fifo_next1<54> ,
         \fifo_next1<53> , \fifo_next1<52> , \fifo_next1<51> ,
         \fifo_next1<50> , \fifo_next1<49> , \fifo_next1<48> ,
         \fifo_next1<47> , \fifo_next1<46> , \fifo_next1<45> ,
         \fifo_next1<44> , \fifo_next1<43> , \fifo_next1<42> ,
         \fifo_next1<41> , \fifo_next1<40> , \fifo_next1<39> ,
         \fifo_next1<38> , \fifo_next1<37> , \fifo_next1<36> ,
         \fifo_next1<35> , \fifo_next1<34> , \fifo_next1<33> ,
         \fifo_next1<32> , \fifo_next1<31> , \fifo_next1<30> ,
         \fifo_next1<29> , \fifo_next1<28> , \fifo_next1<27> ,
         \fifo_next1<26> , \fifo_next1<25> , \fifo_next1<24> ,
         \fifo_next1<23> , \fifo_next1<22> , \fifo_next1<21> ,
         \fifo_next1<20> , \fifo_next1<19> , \fifo_next1<18> ,
         \fifo_next1<17> , \fifo_next1<16> , \fifo_next1<15> ,
         \fifo_next1<14> , \fifo_next1<13> , \fifo_next1<12> ,
         \fifo_next1<11> , \fifo_next1<10> , \fifo_next1<9> , \fifo_next1<8> ,
         \fifo_next1<7> , \fifo_next1<6> , \fifo_next1<5> , \fifo_next1<4> ,
         \fifo_next1<3> , \fifo_next1<2> , \fifo_next1<1> , \fifo_next1<0> ,
         \fifo2<63> , \fifo2<62> , \fifo2<61> , \fifo2<60> , \fifo2<59> ,
         \fifo2<58> , \fifo2<57> , \fifo2<56> , \fifo2<55> , \fifo2<54> ,
         \fifo2<53> , \fifo2<52> , \fifo2<51> , \fifo2<50> , \fifo2<49> ,
         \fifo2<48> , \fifo2<47> , \fifo2<46> , \fifo2<45> , \fifo2<44> ,
         \fifo2<43> , \fifo2<42> , \fifo2<41> , \fifo2<40> , \fifo2<39> ,
         \fifo2<38> , \fifo2<37> , \fifo2<36> , \fifo2<35> , \fifo2<34> ,
         \fifo2<33> , \fifo2<32> , \fifo2<31> , \fifo2<30> , \fifo2<29> ,
         \fifo2<28> , \fifo2<27> , \fifo2<26> , \fifo2<25> , \fifo2<24> ,
         \fifo2<23> , \fifo2<22> , \fifo2<21> , \fifo2<20> , \fifo2<19> ,
         \fifo2<18> , \fifo2<17> , \fifo2<16> , \fifo2<15> , \fifo2<14> ,
         \fifo2<13> , \fifo2<12> , \fifo2<11> , \fifo2<10> , \fifo2<9> ,
         \fifo2<8> , \fifo2<7> , \fifo2<6> , \fifo2<5> , \fifo2<4> ,
         \fifo2<3> , \fifo2<2> , \fifo2<1> , \fifo2<0> , \fifo_next2<63> ,
         \fifo_next2<62> , \fifo_next2<61> , \fifo_next2<60> ,
         \fifo_next2<59> , \fifo_next2<58> , \fifo_next2<57> ,
         \fifo_next2<56> , \fifo_next2<55> , \fifo_next2<54> ,
         \fifo_next2<53> , \fifo_next2<52> , \fifo_next2<51> ,
         \fifo_next2<50> , \fifo_next2<49> , \fifo_next2<48> ,
         \fifo_next2<47> , \fifo_next2<46> , \fifo_next2<45> ,
         \fifo_next2<44> , \fifo_next2<43> , \fifo_next2<42> ,
         \fifo_next2<41> , \fifo_next2<40> , \fifo_next2<39> ,
         \fifo_next2<38> , \fifo_next2<37> , \fifo_next2<36> ,
         \fifo_next2<35> , \fifo_next2<34> , \fifo_next2<33> ,
         \fifo_next2<32> , \fifo_next2<31> , \fifo_next2<30> ,
         \fifo_next2<29> , \fifo_next2<28> , \fifo_next2<27> ,
         \fifo_next2<26> , \fifo_next2<25> , \fifo_next2<24> ,
         \fifo_next2<23> , \fifo_next2<22> , \fifo_next2<21> ,
         \fifo_next2<20> , \fifo_next2<19> , \fifo_next2<18> ,
         \fifo_next2<17> , \fifo_next2<16> , \fifo_next2<15> ,
         \fifo_next2<14> , \fifo_next2<13> , \fifo_next2<12> ,
         \fifo_next2<11> , \fifo_next2<10> , \fifo_next2<9> , \fifo_next2<8> ,
         \fifo_next2<7> , \fifo_next2<6> , \fifo_next2<5> , \fifo_next2<4> ,
         \fifo_next2<3> , \fifo_next2<2> , \fifo_next2<1> , \fifo_next2<0> ,
         \fifo3<63> , \fifo3<62> , \fifo3<61> , \fifo3<60> , \fifo3<59> ,
         \fifo3<58> , \fifo3<57> , \fifo3<56> , \fifo3<55> , \fifo3<54> ,
         \fifo3<53> , \fifo3<52> , \fifo3<51> , \fifo3<50> , \fifo3<49> ,
         \fifo3<48> , \fifo3<47> , \fifo3<46> , \fifo3<45> , \fifo3<44> ,
         \fifo3<43> , \fifo3<42> , \fifo3<41> , \fifo3<40> , \fifo3<39> ,
         \fifo3<38> , \fifo3<37> , \fifo3<36> , \fifo3<35> , \fifo3<34> ,
         \fifo3<33> , \fifo3<32> , \fifo3<31> , \fifo3<30> , \fifo3<29> ,
         \fifo3<28> , \fifo3<27> , \fifo3<26> , \fifo3<25> , \fifo3<24> ,
         \fifo3<23> , \fifo3<22> , \fifo3<21> , \fifo3<20> , \fifo3<19> ,
         \fifo3<18> , \fifo3<17> , \fifo3<16> , \fifo3<15> , \fifo3<14> ,
         \fifo3<13> , \fifo3<12> , \fifo3<11> , \fifo3<10> , \fifo3<9> ,
         \fifo3<8> , \fifo3<7> , \fifo3<6> , \fifo3<5> , \fifo3<4> ,
         \fifo3<3> , \fifo3<2> , \fifo3<1> , \fifo3<0> , \fifo_next3<63> ,
         \fifo_next3<62> , \fifo_next3<61> , \fifo_next3<60> ,
         \fifo_next3<59> , \fifo_next3<58> , \fifo_next3<57> ,
         \fifo_next3<56> , \fifo_next3<55> , \fifo_next3<54> ,
         \fifo_next3<53> , \fifo_next3<52> , \fifo_next3<51> ,
         \fifo_next3<50> , \fifo_next3<49> , \fifo_next3<48> ,
         \fifo_next3<47> , \fifo_next3<46> , \fifo_next3<45> ,
         \fifo_next3<44> , \fifo_next3<43> , \fifo_next3<42> ,
         \fifo_next3<41> , \fifo_next3<40> , \fifo_next3<39> ,
         \fifo_next3<38> , \fifo_next3<37> , \fifo_next3<36> ,
         \fifo_next3<35> , \fifo_next3<34> , \fifo_next3<33> ,
         \fifo_next3<32> , \fifo_next3<31> , \fifo_next3<30> ,
         \fifo_next3<29> , \fifo_next3<28> , \fifo_next3<27> ,
         \fifo_next3<26> , \fifo_next3<25> , \fifo_next3<24> ,
         \fifo_next3<23> , \fifo_next3<22> , \fifo_next3<21> ,
         \fifo_next3<20> , \fifo_next3<19> , \fifo_next3<18> ,
         \fifo_next3<17> , \fifo_next3<16> , \fifo_next3<15> ,
         \fifo_next3<14> , \fifo_next3<13> , \fifo_next3<12> ,
         \fifo_next3<11> , \fifo_next3<10> , \fifo_next3<9> , \fifo_next3<8> ,
         \fifo_next3<7> , \fifo_next3<6> , \fifo_next3<5> , \fifo_next3<4> ,
         \fifo_next3<3> , \fifo_next3<2> , \fifo_next3<1> , \fifo_next3<0> ,
         \readstate<1> , \readstate<0> , \readstate_plus1<1> ,
         \readstate_plus1<0> , \writestate<1> , \writestate<0> ,
         \writestate_plus1<1> , \writestate_plus1<0> , \rwcounter<3> ,
         \rwcounter<2> , \rwcounter<1> , \rwcounter<0> , \readstate_next<1> ,
         \readstate_next<0> , n10, n12, n16, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667;

  AOI22X1 U17 ( .A(\writestate<1> ), .B(n152), .C(\writestate_plus1<1> ), .D(
        n306), .Y(n10) );
  AOI22X1 U18 ( .A(\writestate<0> ), .B(n152), .C(\writestate_plus1<0> ), .D(
        n306), .Y(n12) );
  OAI21X1 U20 ( .A(data_out_valid), .B(n666), .C(n156), .Y(\readstate_next<1> ) );
  OAI21X1 U22 ( .A(data_out_valid), .B(n665), .C(n154), .Y(\readstate_next<0> ) );
  NOR3X1 U26 ( .A(\rwcounter<0> ), .B(\rwcounter<3> ), .C(\rwcounter<1> ), .Y(
        n16) );
  NAND2X1 U27 ( .A(n284), .B(n220), .Y(\data_out<9> ) );
  AOI22X1 U28 ( .A(\fifo3<9> ), .B(n656), .C(\fifo2<9> ), .D(n21), .Y(n19) );
  AOI22X1 U29 ( .A(\fifo1<9> ), .B(n22), .C(\fifo0<9> ), .D(n645), .Y(n18) );
  NAND2X1 U30 ( .A(n283), .B(n219), .Y(\data_out<8> ) );
  AOI22X1 U31 ( .A(\fifo3<8> ), .B(n656), .C(\fifo2<8> ), .D(n21), .Y(n25) );
  AOI22X1 U32 ( .A(\fifo1<8> ), .B(n22), .C(\fifo0<8> ), .D(n23), .Y(n24) );
  NAND2X1 U33 ( .A(n282), .B(n218), .Y(\data_out<7> ) );
  AOI22X1 U34 ( .A(\fifo3<7> ), .B(n656), .C(\fifo2<7> ), .D(n21), .Y(n27) );
  AOI22X1 U35 ( .A(\fifo1<7> ), .B(n22), .C(\fifo0<7> ), .D(n645), .Y(n26) );
  NAND2X1 U36 ( .A(n281), .B(n217), .Y(\data_out<6> ) );
  AOI22X1 U37 ( .A(\fifo3<6> ), .B(n656), .C(\fifo2<6> ), .D(n21), .Y(n29) );
  AOI22X1 U38 ( .A(\fifo1<6> ), .B(n22), .C(\fifo0<6> ), .D(n23), .Y(n28) );
  NAND2X1 U39 ( .A(n280), .B(n216), .Y(\data_out<63> ) );
  AOI22X1 U40 ( .A(\fifo3<63> ), .B(n656), .C(\fifo2<63> ), .D(n21), .Y(n31)
         );
  AOI22X1 U41 ( .A(\fifo1<63> ), .B(n22), .C(\fifo0<63> ), .D(n645), .Y(n30)
         );
  NAND2X1 U42 ( .A(n279), .B(n215), .Y(\data_out<62> ) );
  AOI22X1 U43 ( .A(\fifo3<62> ), .B(n656), .C(\fifo2<62> ), .D(n21), .Y(n33)
         );
  AOI22X1 U44 ( .A(\fifo1<62> ), .B(n22), .C(\fifo0<62> ), .D(n23), .Y(n32) );
  NAND2X1 U45 ( .A(n278), .B(n214), .Y(\data_out<61> ) );
  AOI22X1 U46 ( .A(\fifo3<61> ), .B(n656), .C(\fifo2<61> ), .D(n21), .Y(n35)
         );
  AOI22X1 U47 ( .A(\fifo1<61> ), .B(n22), .C(\fifo0<61> ), .D(n645), .Y(n34)
         );
  NAND2X1 U48 ( .A(n277), .B(n213), .Y(\data_out<60> ) );
  AOI22X1 U49 ( .A(\fifo3<60> ), .B(n656), .C(\fifo2<60> ), .D(n21), .Y(n37)
         );
  AOI22X1 U50 ( .A(\fifo1<60> ), .B(n22), .C(\fifo0<60> ), .D(n645), .Y(n36)
         );
  NAND2X1 U51 ( .A(n276), .B(n212), .Y(\data_out<5> ) );
  AOI22X1 U52 ( .A(\fifo3<5> ), .B(n656), .C(\fifo2<5> ), .D(n21), .Y(n39) );
  AOI22X1 U53 ( .A(\fifo1<5> ), .B(n22), .C(\fifo0<5> ), .D(n645), .Y(n38) );
  NAND2X1 U54 ( .A(n275), .B(n211), .Y(\data_out<59> ) );
  AOI22X1 U55 ( .A(\fifo3<59> ), .B(n656), .C(\fifo2<59> ), .D(n21), .Y(n41)
         );
  AOI22X1 U56 ( .A(\fifo1<59> ), .B(n22), .C(\fifo0<59> ), .D(n645), .Y(n40)
         );
  NAND2X1 U57 ( .A(n274), .B(n210), .Y(\data_out<58> ) );
  AOI22X1 U58 ( .A(\fifo3<58> ), .B(n656), .C(\fifo2<58> ), .D(n21), .Y(n43)
         );
  AOI22X1 U59 ( .A(\fifo1<58> ), .B(n22), .C(\fifo0<58> ), .D(n645), .Y(n42)
         );
  NAND2X1 U60 ( .A(n273), .B(n209), .Y(\data_out<57> ) );
  AOI22X1 U61 ( .A(\fifo3<57> ), .B(n656), .C(\fifo2<57> ), .D(n21), .Y(n45)
         );
  AOI22X1 U62 ( .A(\fifo1<57> ), .B(n22), .C(\fifo0<57> ), .D(n645), .Y(n44)
         );
  NAND2X1 U63 ( .A(n272), .B(n208), .Y(\data_out<56> ) );
  AOI22X1 U64 ( .A(\fifo3<56> ), .B(n656), .C(\fifo2<56> ), .D(n21), .Y(n47)
         );
  AOI22X1 U65 ( .A(\fifo1<56> ), .B(n22), .C(\fifo0<56> ), .D(n23), .Y(n46) );
  NAND2X1 U66 ( .A(n271), .B(n207), .Y(\data_out<55> ) );
  AOI22X1 U67 ( .A(\fifo3<55> ), .B(n20), .C(\fifo2<55> ), .D(n21), .Y(n49) );
  AOI22X1 U68 ( .A(\fifo1<55> ), .B(n648), .C(\fifo0<55> ), .D(n23), .Y(n48)
         );
  NAND2X1 U69 ( .A(n270), .B(n206), .Y(\data_out<54> ) );
  AOI22X1 U70 ( .A(\fifo3<54> ), .B(n20), .C(\fifo2<54> ), .D(n21), .Y(n51) );
  AOI22X1 U71 ( .A(\fifo1<54> ), .B(n648), .C(\fifo0<54> ), .D(n23), .Y(n50)
         );
  NAND2X1 U72 ( .A(n269), .B(n205), .Y(\data_out<53> ) );
  AOI22X1 U73 ( .A(\fifo3<53> ), .B(n20), .C(\fifo2<53> ), .D(n21), .Y(n53) );
  AOI22X1 U74 ( .A(\fifo1<53> ), .B(n648), .C(\fifo0<53> ), .D(n23), .Y(n52)
         );
  NAND2X1 U75 ( .A(n268), .B(n204), .Y(\data_out<52> ) );
  AOI22X1 U76 ( .A(\fifo3<52> ), .B(n20), .C(\fifo2<52> ), .D(n21), .Y(n55) );
  AOI22X1 U77 ( .A(\fifo1<52> ), .B(n648), .C(\fifo0<52> ), .D(n23), .Y(n54)
         );
  NAND2X1 U78 ( .A(n267), .B(n203), .Y(\data_out<51> ) );
  AOI22X1 U79 ( .A(\fifo3<51> ), .B(n20), .C(\fifo2<51> ), .D(n21), .Y(n57) );
  AOI22X1 U80 ( .A(\fifo1<51> ), .B(n648), .C(\fifo0<51> ), .D(n23), .Y(n56)
         );
  NAND2X1 U81 ( .A(n266), .B(n202), .Y(\data_out<50> ) );
  AOI22X1 U82 ( .A(\fifo3<50> ), .B(n20), .C(\fifo2<50> ), .D(n21), .Y(n59) );
  AOI22X1 U83 ( .A(\fifo1<50> ), .B(n648), .C(\fifo0<50> ), .D(n23), .Y(n58)
         );
  NAND2X1 U84 ( .A(n265), .B(n201), .Y(\data_out<4> ) );
  AOI22X1 U85 ( .A(\fifo3<4> ), .B(n20), .C(\fifo2<4> ), .D(n21), .Y(n61) );
  AOI22X1 U86 ( .A(\fifo1<4> ), .B(n648), .C(\fifo0<4> ), .D(n23), .Y(n60) );
  NAND2X1 U87 ( .A(n264), .B(n200), .Y(\data_out<49> ) );
  AOI22X1 U88 ( .A(\fifo3<49> ), .B(n20), .C(\fifo2<49> ), .D(n21), .Y(n63) );
  AOI22X1 U89 ( .A(\fifo1<49> ), .B(n648), .C(\fifo0<49> ), .D(n23), .Y(n62)
         );
  NAND2X1 U90 ( .A(n263), .B(n199), .Y(\data_out<48> ) );
  AOI22X1 U91 ( .A(\fifo3<48> ), .B(n20), .C(\fifo2<48> ), .D(n21), .Y(n65) );
  AOI22X1 U92 ( .A(\fifo1<48> ), .B(n648), .C(\fifo0<48> ), .D(n23), .Y(n64)
         );
  NAND2X1 U93 ( .A(n262), .B(n198), .Y(\data_out<47> ) );
  AOI22X1 U94 ( .A(\fifo3<47> ), .B(n20), .C(\fifo2<47> ), .D(n21), .Y(n67) );
  AOI22X1 U95 ( .A(\fifo1<47> ), .B(n648), .C(\fifo0<47> ), .D(n23), .Y(n66)
         );
  NAND2X1 U96 ( .A(n261), .B(n197), .Y(\data_out<46> ) );
  AOI22X1 U97 ( .A(\fifo3<46> ), .B(n20), .C(\fifo2<46> ), .D(n21), .Y(n69) );
  AOI22X1 U98 ( .A(\fifo1<46> ), .B(n648), .C(\fifo0<46> ), .D(n23), .Y(n68)
         );
  NAND2X1 U99 ( .A(n260), .B(n196), .Y(\data_out<45> ) );
  AOI22X1 U100 ( .A(\fifo3<45> ), .B(n20), .C(\fifo2<45> ), .D(n652), .Y(n71)
         );
  AOI22X1 U101 ( .A(\fifo1<45> ), .B(n648), .C(\fifo0<45> ), .D(n645), .Y(n70)
         );
  NAND2X1 U102 ( .A(n259), .B(n195), .Y(\data_out<44> ) );
  AOI22X1 U103 ( .A(\fifo3<44> ), .B(n20), .C(\fifo2<44> ), .D(n652), .Y(n73)
         );
  AOI22X1 U104 ( .A(\fifo1<44> ), .B(n648), .C(\fifo0<44> ), .D(n645), .Y(n72)
         );
  NAND2X1 U105 ( .A(n258), .B(n194), .Y(\data_out<43> ) );
  AOI22X1 U106 ( .A(\fifo3<43> ), .B(n20), .C(\fifo2<43> ), .D(n652), .Y(n75)
         );
  AOI22X1 U107 ( .A(\fifo1<43> ), .B(n649), .C(\fifo0<43> ), .D(n645), .Y(n74)
         );
  NAND2X1 U108 ( .A(n257), .B(n193), .Y(\data_out<42> ) );
  AOI22X1 U109 ( .A(\fifo3<42> ), .B(n20), .C(\fifo2<42> ), .D(n652), .Y(n77)
         );
  AOI22X1 U110 ( .A(\fifo1<42> ), .B(n649), .C(\fifo0<42> ), .D(n645), .Y(n76)
         );
  NAND2X1 U111 ( .A(n256), .B(n192), .Y(\data_out<41> ) );
  AOI22X1 U112 ( .A(\fifo3<41> ), .B(n20), .C(\fifo2<41> ), .D(n652), .Y(n79)
         );
  AOI22X1 U113 ( .A(\fifo1<41> ), .B(n649), .C(\fifo0<41> ), .D(n645), .Y(n78)
         );
  NAND2X1 U114 ( .A(n255), .B(n191), .Y(\data_out<40> ) );
  AOI22X1 U115 ( .A(\fifo3<40> ), .B(n20), .C(\fifo2<40> ), .D(n652), .Y(n81)
         );
  AOI22X1 U116 ( .A(\fifo1<40> ), .B(n649), .C(\fifo0<40> ), .D(n645), .Y(n80)
         );
  NAND2X1 U117 ( .A(n254), .B(n190), .Y(\data_out<3> ) );
  AOI22X1 U118 ( .A(\fifo3<3> ), .B(n20), .C(\fifo2<3> ), .D(n652), .Y(n83) );
  AOI22X1 U119 ( .A(\fifo1<3> ), .B(n649), .C(\fifo0<3> ), .D(n645), .Y(n82)
         );
  NAND2X1 U120 ( .A(n253), .B(n189), .Y(\data_out<39> ) );
  AOI22X1 U121 ( .A(\fifo3<39> ), .B(n20), .C(\fifo2<39> ), .D(n652), .Y(n85)
         );
  AOI22X1 U122 ( .A(\fifo1<39> ), .B(n649), .C(\fifo0<39> ), .D(n645), .Y(n84)
         );
  NAND2X1 U123 ( .A(n252), .B(n188), .Y(\data_out<38> ) );
  AOI22X1 U124 ( .A(\fifo3<38> ), .B(n20), .C(\fifo2<38> ), .D(n652), .Y(n87)
         );
  AOI22X1 U125 ( .A(\fifo1<38> ), .B(n649), .C(\fifo0<38> ), .D(n645), .Y(n86)
         );
  NAND2X1 U126 ( .A(n251), .B(n187), .Y(\data_out<37> ) );
  AOI22X1 U127 ( .A(\fifo3<37> ), .B(n20), .C(\fifo2<37> ), .D(n652), .Y(n89)
         );
  AOI22X1 U128 ( .A(\fifo1<37> ), .B(n649), .C(\fifo0<37> ), .D(n645), .Y(n88)
         );
  NAND2X1 U129 ( .A(n250), .B(n186), .Y(\data_out<36> ) );
  AOI22X1 U130 ( .A(\fifo3<36> ), .B(n20), .C(\fifo2<36> ), .D(n652), .Y(n91)
         );
  AOI22X1 U131 ( .A(\fifo1<36> ), .B(n649), .C(\fifo0<36> ), .D(n645), .Y(n90)
         );
  NAND2X1 U132 ( .A(n249), .B(n185), .Y(\data_out<35> ) );
  AOI22X1 U133 ( .A(\fifo3<35> ), .B(n20), .C(\fifo2<35> ), .D(n652), .Y(n93)
         );
  AOI22X1 U134 ( .A(\fifo1<35> ), .B(n649), .C(\fifo0<35> ), .D(n645), .Y(n92)
         );
  NAND2X1 U135 ( .A(n248), .B(n184), .Y(\data_out<34> ) );
  AOI22X1 U136 ( .A(\fifo3<34> ), .B(n20), .C(\fifo2<34> ), .D(n653), .Y(n95)
         );
  AOI22X1 U137 ( .A(\fifo1<34> ), .B(n649), .C(\fifo0<34> ), .D(n23), .Y(n94)
         );
  NAND2X1 U138 ( .A(n247), .B(n183), .Y(\data_out<33> ) );
  AOI22X1 U139 ( .A(\fifo3<33> ), .B(n20), .C(\fifo2<33> ), .D(n653), .Y(n97)
         );
  AOI22X1 U140 ( .A(\fifo1<33> ), .B(n649), .C(\fifo0<33> ), .D(n23), .Y(n96)
         );
  NAND2X1 U141 ( .A(n246), .B(n182), .Y(\data_out<32> ) );
  AOI22X1 U142 ( .A(\fifo3<32> ), .B(n20), .C(\fifo2<32> ), .D(n653), .Y(n99)
         );
  AOI22X1 U143 ( .A(\fifo1<32> ), .B(n649), .C(\fifo0<32> ), .D(n23), .Y(n98)
         );
  NAND2X1 U144 ( .A(n245), .B(n181), .Y(\data_out<31> ) );
  AOI22X1 U145 ( .A(\fifo3<31> ), .B(n657), .C(\fifo2<31> ), .D(n653), .Y(n101) );
  AOI22X1 U146 ( .A(\fifo1<31> ), .B(n650), .C(\fifo0<31> ), .D(n23), .Y(n100)
         );
  NAND2X1 U147 ( .A(n244), .B(n180), .Y(\data_out<30> ) );
  AOI22X1 U148 ( .A(\fifo3<30> ), .B(n657), .C(\fifo2<30> ), .D(n653), .Y(n103) );
  AOI22X1 U149 ( .A(\fifo1<30> ), .B(n650), .C(\fifo0<30> ), .D(n23), .Y(n102)
         );
  NAND2X1 U150 ( .A(n243), .B(n179), .Y(\data_out<2> ) );
  AOI22X1 U151 ( .A(\fifo3<2> ), .B(n657), .C(\fifo2<2> ), .D(n653), .Y(n105)
         );
  AOI22X1 U152 ( .A(\fifo1<2> ), .B(n650), .C(\fifo0<2> ), .D(n23), .Y(n104)
         );
  NAND2X1 U153 ( .A(n242), .B(n178), .Y(\data_out<29> ) );
  AOI22X1 U154 ( .A(\fifo3<29> ), .B(n657), .C(\fifo2<29> ), .D(n653), .Y(n107) );
  AOI22X1 U155 ( .A(\fifo1<29> ), .B(n650), .C(\fifo0<29> ), .D(n646), .Y(n106) );
  NAND2X1 U156 ( .A(n241), .B(n177), .Y(\data_out<28> ) );
  AOI22X1 U157 ( .A(\fifo3<28> ), .B(n657), .C(\fifo2<28> ), .D(n653), .Y(n109) );
  AOI22X1 U158 ( .A(\fifo1<28> ), .B(n650), .C(\fifo0<28> ), .D(n646), .Y(n108) );
  NAND2X1 U159 ( .A(n240), .B(n176), .Y(\data_out<27> ) );
  AOI22X1 U160 ( .A(\fifo3<27> ), .B(n657), .C(\fifo2<27> ), .D(n653), .Y(n111) );
  AOI22X1 U161 ( .A(\fifo1<27> ), .B(n650), .C(\fifo0<27> ), .D(n646), .Y(n110) );
  NAND2X1 U162 ( .A(n239), .B(n175), .Y(\data_out<26> ) );
  AOI22X1 U163 ( .A(\fifo3<26> ), .B(n657), .C(\fifo2<26> ), .D(n653), .Y(n113) );
  AOI22X1 U164 ( .A(\fifo1<26> ), .B(n650), .C(\fifo0<26> ), .D(n646), .Y(n112) );
  NAND2X1 U165 ( .A(n238), .B(n174), .Y(\data_out<25> ) );
  AOI22X1 U166 ( .A(\fifo3<25> ), .B(n657), .C(\fifo2<25> ), .D(n653), .Y(n115) );
  AOI22X1 U167 ( .A(\fifo1<25> ), .B(n650), .C(\fifo0<25> ), .D(n646), .Y(n114) );
  NAND2X1 U168 ( .A(n237), .B(n173), .Y(\data_out<24> ) );
  AOI22X1 U169 ( .A(\fifo3<24> ), .B(n657), .C(\fifo2<24> ), .D(n653), .Y(n117) );
  AOI22X1 U170 ( .A(\fifo1<24> ), .B(n650), .C(\fifo0<24> ), .D(n646), .Y(n116) );
  NAND2X1 U171 ( .A(n236), .B(n172), .Y(\data_out<23> ) );
  AOI22X1 U172 ( .A(\fifo3<23> ), .B(n657), .C(\fifo2<23> ), .D(n654), .Y(n119) );
  AOI22X1 U173 ( .A(\fifo1<23> ), .B(n650), .C(\fifo0<23> ), .D(n646), .Y(n118) );
  NAND2X1 U174 ( .A(n235), .B(n171), .Y(\data_out<22> ) );
  AOI22X1 U175 ( .A(\fifo3<22> ), .B(n657), .C(\fifo2<22> ), .D(n654), .Y(n121) );
  AOI22X1 U176 ( .A(\fifo1<22> ), .B(n650), .C(\fifo0<22> ), .D(n646), .Y(n120) );
  NAND2X1 U177 ( .A(n234), .B(n170), .Y(\data_out<21> ) );
  AOI22X1 U178 ( .A(\fifo3<21> ), .B(n657), .C(\fifo2<21> ), .D(n654), .Y(n123) );
  AOI22X1 U179 ( .A(\fifo1<21> ), .B(n650), .C(\fifo0<21> ), .D(n646), .Y(n122) );
  NAND2X1 U180 ( .A(n233), .B(n169), .Y(\data_out<20> ) );
  AOI22X1 U181 ( .A(\fifo3<20> ), .B(n657), .C(\fifo2<20> ), .D(n654), .Y(n125) );
  AOI22X1 U182 ( .A(\fifo1<20> ), .B(n650), .C(\fifo0<20> ), .D(n646), .Y(n124) );
  NAND2X1 U183 ( .A(n232), .B(n168), .Y(\data_out<1> ) );
  AOI22X1 U184 ( .A(\fifo3<1> ), .B(n20), .C(\fifo2<1> ), .D(n654), .Y(n127)
         );
  AOI22X1 U185 ( .A(\fifo1<1> ), .B(n22), .C(\fifo0<1> ), .D(n646), .Y(n126)
         );
  NAND2X1 U186 ( .A(n231), .B(n167), .Y(\data_out<19> ) );
  AOI22X1 U187 ( .A(\fifo3<19> ), .B(n20), .C(\fifo2<19> ), .D(n654), .Y(n129)
         );
  AOI22X1 U188 ( .A(\fifo1<19> ), .B(n22), .C(\fifo0<19> ), .D(n646), .Y(n128)
         );
  NAND2X1 U189 ( .A(n230), .B(n166), .Y(\data_out<18> ) );
  AOI22X1 U190 ( .A(\fifo3<18> ), .B(n20), .C(\fifo2<18> ), .D(n654), .Y(n131)
         );
  AOI22X1 U191 ( .A(\fifo1<18> ), .B(n22), .C(\fifo0<18> ), .D(n646), .Y(n130)
         );
  NAND2X1 U192 ( .A(n229), .B(n165), .Y(\data_out<17> ) );
  AOI22X1 U193 ( .A(\fifo3<17> ), .B(n20), .C(\fifo2<17> ), .D(n654), .Y(n133)
         );
  AOI22X1 U194 ( .A(\fifo1<17> ), .B(n22), .C(\fifo0<17> ), .D(n646), .Y(n132)
         );
  NAND2X1 U195 ( .A(n228), .B(n164), .Y(\data_out<16> ) );
  AOI22X1 U196 ( .A(\fifo3<16> ), .B(n20), .C(\fifo2<16> ), .D(n654), .Y(n135)
         );
  AOI22X1 U197 ( .A(\fifo1<16> ), .B(n22), .C(\fifo0<16> ), .D(n646), .Y(n134)
         );
  NAND2X1 U198 ( .A(n227), .B(n163), .Y(\data_out<15> ) );
  AOI22X1 U199 ( .A(\fifo3<15> ), .B(n20), .C(\fifo2<15> ), .D(n654), .Y(n137)
         );
  AOI22X1 U200 ( .A(\fifo1<15> ), .B(n22), .C(\fifo0<15> ), .D(n646), .Y(n136)
         );
  NAND2X1 U201 ( .A(n226), .B(n162), .Y(\data_out<14> ) );
  AOI22X1 U202 ( .A(\fifo3<14> ), .B(n20), .C(\fifo2<14> ), .D(n654), .Y(n139)
         );
  AOI22X1 U203 ( .A(\fifo1<14> ), .B(n22), .C(\fifo0<14> ), .D(n646), .Y(n138)
         );
  NAND2X1 U204 ( .A(n225), .B(n161), .Y(\data_out<13> ) );
  AOI22X1 U205 ( .A(\fifo3<13> ), .B(n20), .C(\fifo2<13> ), .D(n654), .Y(n141)
         );
  AOI22X1 U206 ( .A(\fifo1<13> ), .B(n22), .C(\fifo0<13> ), .D(n646), .Y(n140)
         );
  NAND2X1 U207 ( .A(n224), .B(n160), .Y(\data_out<12> ) );
  AOI22X1 U208 ( .A(\fifo3<12> ), .B(n20), .C(\fifo2<12> ), .D(n21), .Y(n143)
         );
  AOI22X1 U209 ( .A(\fifo1<12> ), .B(n22), .C(\fifo0<12> ), .D(n646), .Y(n142)
         );
  NAND2X1 U210 ( .A(n223), .B(n159), .Y(\data_out<11> ) );
  AOI22X1 U211 ( .A(\fifo3<11> ), .B(n20), .C(\fifo2<11> ), .D(n21), .Y(n145)
         );
  AOI22X1 U212 ( .A(\fifo1<11> ), .B(n22), .C(\fifo0<11> ), .D(n23), .Y(n144)
         );
  NAND2X1 U213 ( .A(n222), .B(n158), .Y(\data_out<10> ) );
  AOI22X1 U214 ( .A(\fifo3<10> ), .B(n20), .C(\fifo2<10> ), .D(n21), .Y(n147)
         );
  AOI22X1 U215 ( .A(\fifo1<10> ), .B(n22), .C(\fifo0<10> ), .D(n646), .Y(n146)
         );
  NAND2X1 U216 ( .A(n221), .B(n157), .Y(\data_out<0> ) );
  AOI22X1 U217 ( .A(\fifo3<0> ), .B(n20), .C(\fifo2<0> ), .D(n21), .Y(n149) );
  AOI22X1 U218 ( .A(\fifo1<0> ), .B(n22), .C(\fifo0<0> ), .D(n23), .Y(n148) );
  dff_200 \reg1[0]  ( .q(\fifo0<0> ), .d(\fifo_next0<0> ), .clk(clk), .rst(
        n661) );
  dff_201 \reg1[1]  ( .q(\fifo0<1> ), .d(\fifo_next0<1> ), .clk(clk), .rst(
        n660) );
  dff_202 \reg1[2]  ( .q(\fifo0<2> ), .d(\fifo_next0<2> ), .clk(clk), .rst(
        n662) );
  dff_203 \reg1[3]  ( .q(\fifo0<3> ), .d(\fifo_next0<3> ), .clk(clk), .rst(
        n662) );
  dff_204 \reg1[4]  ( .q(\fifo0<4> ), .d(\fifo_next0<4> ), .clk(clk), .rst(
        n661) );
  dff_205 \reg1[5]  ( .q(\fifo0<5> ), .d(\fifo_next0<5> ), .clk(clk), .rst(
        n662) );
  dff_206 \reg1[6]  ( .q(\fifo0<6> ), .d(\fifo_next0<6> ), .clk(clk), .rst(
        n661) );
  dff_207 \reg1[7]  ( .q(\fifo0<7> ), .d(\fifo_next0<7> ), .clk(clk), .rst(
        n662) );
  dff_208 \reg1[8]  ( .q(\fifo0<8> ), .d(\fifo_next0<8> ), .clk(clk), .rst(
        n661) );
  dff_209 \reg1[9]  ( .q(\fifo0<9> ), .d(\fifo_next0<9> ), .clk(clk), .rst(
        n662) );
  dff_210 \reg1[10]  ( .q(\fifo0<10> ), .d(\fifo_next0<10> ), .clk(clk), .rst(
        n661) );
  dff_211 \reg1[11]  ( .q(\fifo0<11> ), .d(\fifo_next0<11> ), .clk(clk), .rst(
        n662) );
  dff_212 \reg1[12]  ( .q(\fifo0<12> ), .d(\fifo_next0<12> ), .clk(clk), .rst(
        n661) );
  dff_213 \reg1[13]  ( .q(\fifo0<13> ), .d(\fifo_next0<13> ), .clk(clk), .rst(
        n662) );
  dff_214 \reg1[14]  ( .q(\fifo0<14> ), .d(\fifo_next0<14> ), .clk(clk), .rst(
        n661) );
  dff_215 \reg1[15]  ( .q(\fifo0<15> ), .d(\fifo_next0<15> ), .clk(clk), .rst(
        n662) );
  dff_216 \reg1[16]  ( .q(\fifo0<16> ), .d(\fifo_next0<16> ), .clk(clk), .rst(
        n661) );
  dff_217 \reg1[17]  ( .q(\fifo0<17> ), .d(\fifo_next0<17> ), .clk(clk), .rst(
        n662) );
  dff_218 \reg1[18]  ( .q(\fifo0<18> ), .d(\fifo_next0<18> ), .clk(clk), .rst(
        n661) );
  dff_219 \reg1[19]  ( .q(\fifo0<19> ), .d(\fifo_next0<19> ), .clk(clk), .rst(
        n662) );
  dff_220 \reg1[20]  ( .q(\fifo0<20> ), .d(\fifo_next0<20> ), .clk(clk), .rst(
        n661) );
  dff_221 \reg1[21]  ( .q(\fifo0<21> ), .d(\fifo_next0<21> ), .clk(clk), .rst(
        n662) );
  dff_222 \reg1[22]  ( .q(\fifo0<22> ), .d(\fifo_next0<22> ), .clk(clk), .rst(
        n661) );
  dff_223 \reg1[23]  ( .q(\fifo0<23> ), .d(\fifo_next0<23> ), .clk(clk), .rst(
        n662) );
  dff_224 \reg1[24]  ( .q(\fifo0<24> ), .d(\fifo_next0<24> ), .clk(clk), .rst(
        n661) );
  dff_225 \reg1[25]  ( .q(\fifo0<25> ), .d(\fifo_next0<25> ), .clk(clk), .rst(
        n662) );
  dff_226 \reg1[26]  ( .q(\fifo0<26> ), .d(\fifo_next0<26> ), .clk(clk), .rst(
        n661) );
  dff_227 \reg1[27]  ( .q(\fifo0<27> ), .d(\fifo_next0<27> ), .clk(clk), .rst(
        n662) );
  dff_228 \reg1[28]  ( .q(\fifo0<28> ), .d(\fifo_next0<28> ), .clk(clk), .rst(
        n661) );
  dff_229 \reg1[29]  ( .q(\fifo0<29> ), .d(\fifo_next0<29> ), .clk(clk), .rst(
        n662) );
  dff_230 \reg1[30]  ( .q(\fifo0<30> ), .d(\fifo_next0<30> ), .clk(clk), .rst(
        n661) );
  dff_231 \reg1[31]  ( .q(\fifo0<31> ), .d(\fifo_next0<31> ), .clk(clk), .rst(
        n662) );
  dff_232 \reg1[32]  ( .q(\fifo0<32> ), .d(\fifo_next0<32> ), .clk(clk), .rst(
        n661) );
  dff_233 \reg1[33]  ( .q(\fifo0<33> ), .d(\fifo_next0<33> ), .clk(clk), .rst(
        n662) );
  dff_234 \reg1[34]  ( .q(\fifo0<34> ), .d(\fifo_next0<34> ), .clk(clk), .rst(
        n662) );
  dff_235 \reg1[35]  ( .q(\fifo0<35> ), .d(\fifo_next0<35> ), .clk(clk), .rst(
        n662) );
  dff_236 \reg1[36]  ( .q(\fifo0<36> ), .d(\fifo_next0<36> ), .clk(clk), .rst(
        n662) );
  dff_237 \reg1[37]  ( .q(\fifo0<37> ), .d(\fifo_next0<37> ), .clk(clk), .rst(
        n662) );
  dff_238 \reg1[38]  ( .q(\fifo0<38> ), .d(\fifo_next0<38> ), .clk(clk), .rst(
        n662) );
  dff_239 \reg1[39]  ( .q(\fifo0<39> ), .d(\fifo_next0<39> ), .clk(clk), .rst(
        n662) );
  dff_240 \reg1[40]  ( .q(\fifo0<40> ), .d(\fifo_next0<40> ), .clk(clk), .rst(
        n662) );
  dff_241 \reg1[41]  ( .q(\fifo0<41> ), .d(\fifo_next0<41> ), .clk(clk), .rst(
        n662) );
  dff_242 \reg1[42]  ( .q(\fifo0<42> ), .d(\fifo_next0<42> ), .clk(clk), .rst(
        n662) );
  dff_243 \reg1[43]  ( .q(\fifo0<43> ), .d(\fifo_next0<43> ), .clk(clk), .rst(
        n662) );
  dff_244 \reg1[44]  ( .q(\fifo0<44> ), .d(\fifo_next0<44> ), .clk(clk), .rst(
        n662) );
  dff_245 \reg1[45]  ( .q(\fifo0<45> ), .d(\fifo_next0<45> ), .clk(clk), .rst(
        n662) );
  dff_246 \reg1[46]  ( .q(\fifo0<46> ), .d(\fifo_next0<46> ), .clk(clk), .rst(
        n662) );
  dff_247 \reg1[47]  ( .q(\fifo0<47> ), .d(\fifo_next0<47> ), .clk(clk), .rst(
        n662) );
  dff_248 \reg1[48]  ( .q(\fifo0<48> ), .d(\fifo_next0<48> ), .clk(clk), .rst(
        n662) );
  dff_249 \reg1[49]  ( .q(\fifo0<49> ), .d(\fifo_next0<49> ), .clk(clk), .rst(
        n662) );
  dff_250 \reg1[50]  ( .q(\fifo0<50> ), .d(\fifo_next0<50> ), .clk(clk), .rst(
        n662) );
  dff_251 \reg1[51]  ( .q(\fifo0<51> ), .d(\fifo_next0<51> ), .clk(clk), .rst(
        n662) );
  dff_252 \reg1[52]  ( .q(\fifo0<52> ), .d(\fifo_next0<52> ), .clk(clk), .rst(
        n662) );
  dff_253 \reg1[53]  ( .q(\fifo0<53> ), .d(\fifo_next0<53> ), .clk(clk), .rst(
        n662) );
  dff_254 \reg1[54]  ( .q(\fifo0<54> ), .d(\fifo_next0<54> ), .clk(clk), .rst(
        n662) );
  dff_255 \reg1[55]  ( .q(\fifo0<55> ), .d(\fifo_next0<55> ), .clk(clk), .rst(
        n662) );
  dff_256 \reg1[56]  ( .q(\fifo0<56> ), .d(\fifo_next0<56> ), .clk(clk), .rst(
        n662) );
  dff_257 \reg1[57]  ( .q(\fifo0<57> ), .d(\fifo_next0<57> ), .clk(clk), .rst(
        n662) );
  dff_258 \reg1[58]  ( .q(\fifo0<58> ), .d(\fifo_next0<58> ), .clk(clk), .rst(
        n662) );
  dff_259 \reg1[59]  ( .q(\fifo0<59> ), .d(\fifo_next0<59> ), .clk(clk), .rst(
        n662) );
  dff_260 \reg1[60]  ( .q(\fifo0<60> ), .d(\fifo_next0<60> ), .clk(clk), .rst(
        n662) );
  dff_261 \reg1[61]  ( .q(\fifo0<61> ), .d(\fifo_next0<61> ), .clk(clk), .rst(
        n662) );
  dff_262 \reg1[62]  ( .q(\fifo0<62> ), .d(\fifo_next0<62> ), .clk(clk), .rst(
        n662) );
  dff_263 \reg1[63]  ( .q(\fifo0<63> ), .d(\fifo_next0<63> ), .clk(clk), .rst(
        n662) );
  dff_136 \reg2[0]  ( .q(\fifo1<0> ), .d(\fifo_next1<0> ), .clk(clk), .rst(
        n662) );
  dff_137 \reg2[1]  ( .q(\fifo1<1> ), .d(\fifo_next1<1> ), .clk(clk), .rst(
        n662) );
  dff_138 \reg2[2]  ( .q(\fifo1<2> ), .d(\fifo_next1<2> ), .clk(clk), .rst(
        n662) );
  dff_139 \reg2[3]  ( .q(\fifo1<3> ), .d(\fifo_next1<3> ), .clk(clk), .rst(
        n662) );
  dff_140 \reg2[4]  ( .q(\fifo1<4> ), .d(\fifo_next1<4> ), .clk(clk), .rst(
        n662) );
  dff_141 \reg2[5]  ( .q(\fifo1<5> ), .d(\fifo_next1<5> ), .clk(clk), .rst(
        n662) );
  dff_142 \reg2[6]  ( .q(\fifo1<6> ), .d(\fifo_next1<6> ), .clk(clk), .rst(
        n662) );
  dff_143 \reg2[7]  ( .q(\fifo1<7> ), .d(\fifo_next1<7> ), .clk(clk), .rst(
        n662) );
  dff_144 \reg2[8]  ( .q(\fifo1<8> ), .d(\fifo_next1<8> ), .clk(clk), .rst(
        n662) );
  dff_145 \reg2[9]  ( .q(\fifo1<9> ), .d(\fifo_next1<9> ), .clk(clk), .rst(
        n662) );
  dff_146 \reg2[10]  ( .q(\fifo1<10> ), .d(\fifo_next1<10> ), .clk(clk), .rst(
        n662) );
  dff_147 \reg2[11]  ( .q(\fifo1<11> ), .d(\fifo_next1<11> ), .clk(clk), .rst(
        n662) );
  dff_148 \reg2[12]  ( .q(\fifo1<12> ), .d(\fifo_next1<12> ), .clk(clk), .rst(
        n662) );
  dff_149 \reg2[13]  ( .q(\fifo1<13> ), .d(\fifo_next1<13> ), .clk(clk), .rst(
        n662) );
  dff_150 \reg2[14]  ( .q(\fifo1<14> ), .d(\fifo_next1<14> ), .clk(clk), .rst(
        n662) );
  dff_151 \reg2[15]  ( .q(\fifo1<15> ), .d(\fifo_next1<15> ), .clk(clk), .rst(
        n662) );
  dff_152 \reg2[16]  ( .q(\fifo1<16> ), .d(\fifo_next1<16> ), .clk(clk), .rst(
        n662) );
  dff_153 \reg2[17]  ( .q(\fifo1<17> ), .d(\fifo_next1<17> ), .clk(clk), .rst(
        n662) );
  dff_154 \reg2[18]  ( .q(\fifo1<18> ), .d(\fifo_next1<18> ), .clk(clk), .rst(
        n662) );
  dff_155 \reg2[19]  ( .q(\fifo1<19> ), .d(\fifo_next1<19> ), .clk(clk), .rst(
        n662) );
  dff_156 \reg2[20]  ( .q(\fifo1<20> ), .d(\fifo_next1<20> ), .clk(clk), .rst(
        n662) );
  dff_157 \reg2[21]  ( .q(\fifo1<21> ), .d(\fifo_next1<21> ), .clk(clk), .rst(
        n662) );
  dff_158 \reg2[22]  ( .q(\fifo1<22> ), .d(\fifo_next1<22> ), .clk(clk), .rst(
        n662) );
  dff_159 \reg2[23]  ( .q(\fifo1<23> ), .d(\fifo_next1<23> ), .clk(clk), .rst(
        n662) );
  dff_160 \reg2[24]  ( .q(\fifo1<24> ), .d(\fifo_next1<24> ), .clk(clk), .rst(
        n661) );
  dff_161 \reg2[25]  ( .q(\fifo1<25> ), .d(\fifo_next1<25> ), .clk(clk), .rst(
        n662) );
  dff_162 \reg2[26]  ( .q(\fifo1<26> ), .d(\fifo_next1<26> ), .clk(clk), .rst(
        n662) );
  dff_163 \reg2[27]  ( .q(\fifo1<27> ), .d(\fifo_next1<27> ), .clk(clk), .rst(
        n661) );
  dff_164 \reg2[28]  ( .q(\fifo1<28> ), .d(\fifo_next1<28> ), .clk(clk), .rst(
        n661) );
  dff_165 \reg2[29]  ( .q(\fifo1<29> ), .d(\fifo_next1<29> ), .clk(clk), .rst(
        n662) );
  dff_166 \reg2[30]  ( .q(\fifo1<30> ), .d(\fifo_next1<30> ), .clk(clk), .rst(
        n661) );
  dff_167 \reg2[31]  ( .q(\fifo1<31> ), .d(\fifo_next1<31> ), .clk(clk), .rst(
        n662) );
  dff_168 \reg2[32]  ( .q(\fifo1<32> ), .d(\fifo_next1<32> ), .clk(clk), .rst(
        n662) );
  dff_169 \reg2[33]  ( .q(\fifo1<33> ), .d(\fifo_next1<33> ), .clk(clk), .rst(
        n661) );
  dff_170 \reg2[34]  ( .q(\fifo1<34> ), .d(\fifo_next1<34> ), .clk(clk), .rst(
        n661) );
  dff_171 \reg2[35]  ( .q(\fifo1<35> ), .d(\fifo_next1<35> ), .clk(clk), .rst(
        n662) );
  dff_172 \reg2[36]  ( .q(\fifo1<36> ), .d(\fifo_next1<36> ), .clk(clk), .rst(
        n661) );
  dff_173 \reg2[37]  ( .q(\fifo1<37> ), .d(\fifo_next1<37> ), .clk(clk), .rst(
        n662) );
  dff_174 \reg2[38]  ( .q(\fifo1<38> ), .d(\fifo_next1<38> ), .clk(clk), .rst(
        n662) );
  dff_175 \reg2[39]  ( .q(\fifo1<39> ), .d(\fifo_next1<39> ), .clk(clk), .rst(
        n661) );
  dff_176 \reg2[40]  ( .q(\fifo1<40> ), .d(\fifo_next1<40> ), .clk(clk), .rst(
        n661) );
  dff_177 \reg2[41]  ( .q(\fifo1<41> ), .d(\fifo_next1<41> ), .clk(clk), .rst(
        n662) );
  dff_178 \reg2[42]  ( .q(\fifo1<42> ), .d(\fifo_next1<42> ), .clk(clk), .rst(
        n661) );
  dff_179 \reg2[43]  ( .q(\fifo1<43> ), .d(\fifo_next1<43> ), .clk(clk), .rst(
        n662) );
  dff_180 \reg2[44]  ( .q(\fifo1<44> ), .d(\fifo_next1<44> ), .clk(clk), .rst(
        n662) );
  dff_181 \reg2[45]  ( .q(\fifo1<45> ), .d(\fifo_next1<45> ), .clk(clk), .rst(
        n661) );
  dff_182 \reg2[46]  ( .q(\fifo1<46> ), .d(\fifo_next1<46> ), .clk(clk), .rst(
        n661) );
  dff_183 \reg2[47]  ( .q(\fifo1<47> ), .d(\fifo_next1<47> ), .clk(clk), .rst(
        n662) );
  dff_184 \reg2[48]  ( .q(\fifo1<48> ), .d(\fifo_next1<48> ), .clk(clk), .rst(
        n661) );
  dff_185 \reg2[49]  ( .q(\fifo1<49> ), .d(\fifo_next1<49> ), .clk(clk), .rst(
        n662) );
  dff_186 \reg2[50]  ( .q(\fifo1<50> ), .d(\fifo_next1<50> ), .clk(clk), .rst(
        n662) );
  dff_187 \reg2[51]  ( .q(\fifo1<51> ), .d(\fifo_next1<51> ), .clk(clk), .rst(
        n661) );
  dff_188 \reg2[52]  ( .q(\fifo1<52> ), .d(\fifo_next1<52> ), .clk(clk), .rst(
        n661) );
  dff_189 \reg2[53]  ( .q(\fifo1<53> ), .d(\fifo_next1<53> ), .clk(clk), .rst(
        n662) );
  dff_190 \reg2[54]  ( .q(\fifo1<54> ), .d(\fifo_next1<54> ), .clk(clk), .rst(
        n661) );
  dff_191 \reg2[55]  ( .q(\fifo1<55> ), .d(\fifo_next1<55> ), .clk(clk), .rst(
        n662) );
  dff_192 \reg2[56]  ( .q(\fifo1<56> ), .d(\fifo_next1<56> ), .clk(clk), .rst(
        n662) );
  dff_193 \reg2[57]  ( .q(\fifo1<57> ), .d(\fifo_next1<57> ), .clk(clk), .rst(
        n661) );
  dff_194 \reg2[58]  ( .q(\fifo1<58> ), .d(\fifo_next1<58> ), .clk(clk), .rst(
        n661) );
  dff_195 \reg2[59]  ( .q(\fifo1<59> ), .d(\fifo_next1<59> ), .clk(clk), .rst(
        n662) );
  dff_196 \reg2[60]  ( .q(\fifo1<60> ), .d(\fifo_next1<60> ), .clk(clk), .rst(
        n661) );
  dff_197 \reg2[61]  ( .q(\fifo1<61> ), .d(\fifo_next1<61> ), .clk(clk), .rst(
        n662) );
  dff_198 \reg2[62]  ( .q(\fifo1<62> ), .d(\fifo_next1<62> ), .clk(clk), .rst(
        n662) );
  dff_199 \reg2[63]  ( .q(\fifo1<63> ), .d(\fifo_next1<63> ), .clk(clk), .rst(
        n661) );
  dff_72 \reg3[0]  ( .q(\fifo2<0> ), .d(\fifo_next2<0> ), .clk(clk), .rst(n661) );
  dff_73 \reg3[1]  ( .q(\fifo2<1> ), .d(\fifo_next2<1> ), .clk(clk), .rst(n662) );
  dff_74 \reg3[2]  ( .q(\fifo2<2> ), .d(\fifo_next2<2> ), .clk(clk), .rst(n661) );
  dff_75 \reg3[3]  ( .q(\fifo2<3> ), .d(\fifo_next2<3> ), .clk(clk), .rst(n662) );
  dff_76 \reg3[4]  ( .q(\fifo2<4> ), .d(\fifo_next2<4> ), .clk(clk), .rst(n661) );
  dff_77 \reg3[5]  ( .q(\fifo2<5> ), .d(\fifo_next2<5> ), .clk(clk), .rst(n660) );
  dff_78 \reg3[6]  ( .q(\fifo2<6> ), .d(\fifo_next2<6> ), .clk(clk), .rst(n660) );
  dff_79 \reg3[7]  ( .q(\fifo2<7> ), .d(\fifo_next2<7> ), .clk(clk), .rst(n660) );
  dff_80 \reg3[8]  ( .q(\fifo2<8> ), .d(\fifo_next2<8> ), .clk(clk), .rst(n660) );
  dff_81 \reg3[9]  ( .q(\fifo2<9> ), .d(\fifo_next2<9> ), .clk(clk), .rst(n660) );
  dff_82 \reg3[10]  ( .q(\fifo2<10> ), .d(\fifo_next2<10> ), .clk(clk), .rst(
        n660) );
  dff_83 \reg3[11]  ( .q(\fifo2<11> ), .d(\fifo_next2<11> ), .clk(clk), .rst(
        n660) );
  dff_84 \reg3[12]  ( .q(\fifo2<12> ), .d(\fifo_next2<12> ), .clk(clk), .rst(
        n660) );
  dff_85 \reg3[13]  ( .q(\fifo2<13> ), .d(\fifo_next2<13> ), .clk(clk), .rst(
        n660) );
  dff_86 \reg3[14]  ( .q(\fifo2<14> ), .d(\fifo_next2<14> ), .clk(clk), .rst(
        n660) );
  dff_87 \reg3[15]  ( .q(\fifo2<15> ), .d(\fifo_next2<15> ), .clk(clk), .rst(
        n660) );
  dff_88 \reg3[16]  ( .q(\fifo2<16> ), .d(\fifo_next2<16> ), .clk(clk), .rst(
        n660) );
  dff_89 \reg3[17]  ( .q(\fifo2<17> ), .d(\fifo_next2<17> ), .clk(clk), .rst(
        n660) );
  dff_90 \reg3[18]  ( .q(\fifo2<18> ), .d(\fifo_next2<18> ), .clk(clk), .rst(
        n660) );
  dff_91 \reg3[19]  ( .q(\fifo2<19> ), .d(\fifo_next2<19> ), .clk(clk), .rst(
        n660) );
  dff_92 \reg3[20]  ( .q(\fifo2<20> ), .d(\fifo_next2<20> ), .clk(clk), .rst(
        n660) );
  dff_93 \reg3[21]  ( .q(\fifo2<21> ), .d(\fifo_next2<21> ), .clk(clk), .rst(
        n660) );
  dff_94 \reg3[22]  ( .q(\fifo2<22> ), .d(\fifo_next2<22> ), .clk(clk), .rst(
        n660) );
  dff_95 \reg3[23]  ( .q(\fifo2<23> ), .d(\fifo_next2<23> ), .clk(clk), .rst(
        n660) );
  dff_96 \reg3[24]  ( .q(\fifo2<24> ), .d(\fifo_next2<24> ), .clk(clk), .rst(
        n660) );
  dff_97 \reg3[25]  ( .q(\fifo2<25> ), .d(\fifo_next2<25> ), .clk(clk), .rst(
        n660) );
  dff_98 \reg3[26]  ( .q(\fifo2<26> ), .d(\fifo_next2<26> ), .clk(clk), .rst(
        n660) );
  dff_99 \reg3[27]  ( .q(\fifo2<27> ), .d(\fifo_next2<27> ), .clk(clk), .rst(
        n660) );
  dff_100 \reg3[28]  ( .q(\fifo2<28> ), .d(\fifo_next2<28> ), .clk(clk), .rst(
        n660) );
  dff_101 \reg3[29]  ( .q(\fifo2<29> ), .d(\fifo_next2<29> ), .clk(clk), .rst(
        n660) );
  dff_102 \reg3[30]  ( .q(\fifo2<30> ), .d(\fifo_next2<30> ), .clk(clk), .rst(
        n660) );
  dff_103 \reg3[31]  ( .q(\fifo2<31> ), .d(\fifo_next2<31> ), .clk(clk), .rst(
        n660) );
  dff_104 \reg3[32]  ( .q(\fifo2<32> ), .d(\fifo_next2<32> ), .clk(clk), .rst(
        n660) );
  dff_105 \reg3[33]  ( .q(\fifo2<33> ), .d(\fifo_next2<33> ), .clk(clk), .rst(
        n660) );
  dff_106 \reg3[34]  ( .q(\fifo2<34> ), .d(\fifo_next2<34> ), .clk(clk), .rst(
        n660) );
  dff_107 \reg3[35]  ( .q(\fifo2<35> ), .d(\fifo_next2<35> ), .clk(clk), .rst(
        n660) );
  dff_108 \reg3[36]  ( .q(\fifo2<36> ), .d(\fifo_next2<36> ), .clk(clk), .rst(
        n660) );
  dff_109 \reg3[37]  ( .q(\fifo2<37> ), .d(\fifo_next2<37> ), .clk(clk), .rst(
        n660) );
  dff_110 \reg3[38]  ( .q(\fifo2<38> ), .d(\fifo_next2<38> ), .clk(clk), .rst(
        n660) );
  dff_111 \reg3[39]  ( .q(\fifo2<39> ), .d(\fifo_next2<39> ), .clk(clk), .rst(
        n660) );
  dff_112 \reg3[40]  ( .q(\fifo2<40> ), .d(\fifo_next2<40> ), .clk(clk), .rst(
        n660) );
  dff_113 \reg3[41]  ( .q(\fifo2<41> ), .d(\fifo_next2<41> ), .clk(clk), .rst(
        n660) );
  dff_114 \reg3[42]  ( .q(\fifo2<42> ), .d(\fifo_next2<42> ), .clk(clk), .rst(
        n660) );
  dff_115 \reg3[43]  ( .q(\fifo2<43> ), .d(\fifo_next2<43> ), .clk(clk), .rst(
        n660) );
  dff_116 \reg3[44]  ( .q(\fifo2<44> ), .d(\fifo_next2<44> ), .clk(clk), .rst(
        n660) );
  dff_117 \reg3[45]  ( .q(\fifo2<45> ), .d(\fifo_next2<45> ), .clk(clk), .rst(
        n660) );
  dff_118 \reg3[46]  ( .q(\fifo2<46> ), .d(\fifo_next2<46> ), .clk(clk), .rst(
        n660) );
  dff_119 \reg3[47]  ( .q(\fifo2<47> ), .d(\fifo_next2<47> ), .clk(clk), .rst(
        n660) );
  dff_120 \reg3[48]  ( .q(\fifo2<48> ), .d(\fifo_next2<48> ), .clk(clk), .rst(
        n660) );
  dff_121 \reg3[49]  ( .q(\fifo2<49> ), .d(\fifo_next2<49> ), .clk(clk), .rst(
        n660) );
  dff_122 \reg3[50]  ( .q(\fifo2<50> ), .d(\fifo_next2<50> ), .clk(clk), .rst(
        n660) );
  dff_123 \reg3[51]  ( .q(\fifo2<51> ), .d(\fifo_next2<51> ), .clk(clk), .rst(
        n660) );
  dff_124 \reg3[52]  ( .q(\fifo2<52> ), .d(\fifo_next2<52> ), .clk(clk), .rst(
        n660) );
  dff_125 \reg3[53]  ( .q(\fifo2<53> ), .d(\fifo_next2<53> ), .clk(clk), .rst(
        n660) );
  dff_126 \reg3[54]  ( .q(\fifo2<54> ), .d(\fifo_next2<54> ), .clk(clk), .rst(
        n661) );
  dff_127 \reg3[55]  ( .q(\fifo2<55> ), .d(\fifo_next2<55> ), .clk(clk), .rst(
        n661) );
  dff_128 \reg3[56]  ( .q(\fifo2<56> ), .d(\fifo_next2<56> ), .clk(clk), .rst(
        n661) );
  dff_129 \reg3[57]  ( .q(\fifo2<57> ), .d(\fifo_next2<57> ), .clk(clk), .rst(
        n661) );
  dff_130 \reg3[58]  ( .q(\fifo2<58> ), .d(\fifo_next2<58> ), .clk(clk), .rst(
        n661) );
  dff_131 \reg3[59]  ( .q(\fifo2<59> ), .d(\fifo_next2<59> ), .clk(clk), .rst(
        n661) );
  dff_132 \reg3[60]  ( .q(\fifo2<60> ), .d(\fifo_next2<60> ), .clk(clk), .rst(
        n661) );
  dff_133 \reg3[61]  ( .q(\fifo2<61> ), .d(\fifo_next2<61> ), .clk(clk), .rst(
        n661) );
  dff_134 \reg3[62]  ( .q(\fifo2<62> ), .d(\fifo_next2<62> ), .clk(clk), .rst(
        n661) );
  dff_135 \reg3[63]  ( .q(\fifo2<63> ), .d(\fifo_next2<63> ), .clk(clk), .rst(
        n661) );
  dff_8 \reg4[0]  ( .q(\fifo3<0> ), .d(\fifo_next3<0> ), .clk(clk), .rst(n661)
         );
  dff_9 \reg4[1]  ( .q(\fifo3<1> ), .d(\fifo_next3<1> ), .clk(clk), .rst(n661)
         );
  dff_10 \reg4[2]  ( .q(\fifo3<2> ), .d(\fifo_next3<2> ), .clk(clk), .rst(n661) );
  dff_11 \reg4[3]  ( .q(\fifo3<3> ), .d(\fifo_next3<3> ), .clk(clk), .rst(n661) );
  dff_12 \reg4[4]  ( .q(\fifo3<4> ), .d(\fifo_next3<4> ), .clk(clk), .rst(n661) );
  dff_13 \reg4[5]  ( .q(\fifo3<5> ), .d(\fifo_next3<5> ), .clk(clk), .rst(n661) );
  dff_14 \reg4[6]  ( .q(\fifo3<6> ), .d(\fifo_next3<6> ), .clk(clk), .rst(n661) );
  dff_15 \reg4[7]  ( .q(\fifo3<7> ), .d(\fifo_next3<7> ), .clk(clk), .rst(n661) );
  dff_16 \reg4[8]  ( .q(\fifo3<8> ), .d(\fifo_next3<8> ), .clk(clk), .rst(n661) );
  dff_17 \reg4[9]  ( .q(\fifo3<9> ), .d(\fifo_next3<9> ), .clk(clk), .rst(n661) );
  dff_18 \reg4[10]  ( .q(\fifo3<10> ), .d(\fifo_next3<10> ), .clk(clk), .rst(
        n661) );
  dff_19 \reg4[11]  ( .q(\fifo3<11> ), .d(\fifo_next3<11> ), .clk(clk), .rst(
        n661) );
  dff_20 \reg4[12]  ( .q(\fifo3<12> ), .d(\fifo_next3<12> ), .clk(clk), .rst(
        n661) );
  dff_21 \reg4[13]  ( .q(\fifo3<13> ), .d(\fifo_next3<13> ), .clk(clk), .rst(
        n661) );
  dff_22 \reg4[14]  ( .q(\fifo3<14> ), .d(\fifo_next3<14> ), .clk(clk), .rst(
        n661) );
  dff_23 \reg4[15]  ( .q(\fifo3<15> ), .d(\fifo_next3<15> ), .clk(clk), .rst(
        n661) );
  dff_24 \reg4[16]  ( .q(\fifo3<16> ), .d(\fifo_next3<16> ), .clk(clk), .rst(
        n661) );
  dff_25 \reg4[17]  ( .q(\fifo3<17> ), .d(\fifo_next3<17> ), .clk(clk), .rst(
        n661) );
  dff_26 \reg4[18]  ( .q(\fifo3<18> ), .d(\fifo_next3<18> ), .clk(clk), .rst(
        n661) );
  dff_27 \reg4[19]  ( .q(\fifo3<19> ), .d(\fifo_next3<19> ), .clk(clk), .rst(
        n661) );
  dff_28 \reg4[20]  ( .q(\fifo3<20> ), .d(\fifo_next3<20> ), .clk(clk), .rst(
        n661) );
  dff_29 \reg4[21]  ( .q(\fifo3<21> ), .d(\fifo_next3<21> ), .clk(clk), .rst(
        n661) );
  dff_30 \reg4[22]  ( .q(\fifo3<22> ), .d(\fifo_next3<22> ), .clk(clk), .rst(
        n661) );
  dff_31 \reg4[23]  ( .q(\fifo3<23> ), .d(\fifo_next3<23> ), .clk(clk), .rst(
        n661) );
  dff_32 \reg4[24]  ( .q(\fifo3<24> ), .d(\fifo_next3<24> ), .clk(clk), .rst(
        n661) );
  dff_33 \reg4[25]  ( .q(\fifo3<25> ), .d(\fifo_next3<25> ), .clk(clk), .rst(
        n661) );
  dff_34 \reg4[26]  ( .q(\fifo3<26> ), .d(\fifo_next3<26> ), .clk(clk), .rst(
        n661) );
  dff_35 \reg4[27]  ( .q(\fifo3<27> ), .d(\fifo_next3<27> ), .clk(clk), .rst(
        n661) );
  dff_36 \reg4[28]  ( .q(\fifo3<28> ), .d(\fifo_next3<28> ), .clk(clk), .rst(
        n661) );
  dff_37 \reg4[29]  ( .q(\fifo3<29> ), .d(\fifo_next3<29> ), .clk(clk), .rst(
        n661) );
  dff_38 \reg4[30]  ( .q(\fifo3<30> ), .d(\fifo_next3<30> ), .clk(clk), .rst(
        n661) );
  dff_39 \reg4[31]  ( .q(\fifo3<31> ), .d(\fifo_next3<31> ), .clk(clk), .rst(
        n661) );
  dff_40 \reg4[32]  ( .q(\fifo3<32> ), .d(\fifo_next3<32> ), .clk(clk), .rst(
        n661) );
  dff_41 \reg4[33]  ( .q(\fifo3<33> ), .d(\fifo_next3<33> ), .clk(clk), .rst(
        n661) );
  dff_42 \reg4[34]  ( .q(\fifo3<34> ), .d(\fifo_next3<34> ), .clk(clk), .rst(
        n661) );
  dff_43 \reg4[35]  ( .q(\fifo3<35> ), .d(\fifo_next3<35> ), .clk(clk), .rst(
        n661) );
  dff_44 \reg4[36]  ( .q(\fifo3<36> ), .d(\fifo_next3<36> ), .clk(clk), .rst(
        n661) );
  dff_45 \reg4[37]  ( .q(\fifo3<37> ), .d(\fifo_next3<37> ), .clk(clk), .rst(
        n661) );
  dff_46 \reg4[38]  ( .q(\fifo3<38> ), .d(\fifo_next3<38> ), .clk(clk), .rst(
        n661) );
  dff_47 \reg4[39]  ( .q(\fifo3<39> ), .d(\fifo_next3<39> ), .clk(clk), .rst(
        n661) );
  dff_48 \reg4[40]  ( .q(\fifo3<40> ), .d(\fifo_next3<40> ), .clk(clk), .rst(
        n661) );
  dff_49 \reg4[41]  ( .q(\fifo3<41> ), .d(\fifo_next3<41> ), .clk(clk), .rst(
        n661) );
  dff_50 \reg4[42]  ( .q(\fifo3<42> ), .d(\fifo_next3<42> ), .clk(clk), .rst(
        n661) );
  dff_51 \reg4[43]  ( .q(\fifo3<43> ), .d(\fifo_next3<43> ), .clk(clk), .rst(
        n661) );
  dff_52 \reg4[44]  ( .q(\fifo3<44> ), .d(\fifo_next3<44> ), .clk(clk), .rst(
        n661) );
  dff_53 \reg4[45]  ( .q(\fifo3<45> ), .d(\fifo_next3<45> ), .clk(clk), .rst(
        n662) );
  dff_54 \reg4[46]  ( .q(\fifo3<46> ), .d(\fifo_next3<46> ), .clk(clk), .rst(
        n661) );
  dff_55 \reg4[47]  ( .q(\fifo3<47> ), .d(\fifo_next3<47> ), .clk(clk), .rst(
        n662) );
  dff_56 \reg4[48]  ( .q(\fifo3<48> ), .d(\fifo_next3<48> ), .clk(clk), .rst(
        n661) );
  dff_57 \reg4[49]  ( .q(\fifo3<49> ), .d(\fifo_next3<49> ), .clk(clk), .rst(
        n662) );
  dff_58 \reg4[50]  ( .q(\fifo3<50> ), .d(\fifo_next3<50> ), .clk(clk), .rst(
        n661) );
  dff_59 \reg4[51]  ( .q(\fifo3<51> ), .d(\fifo_next3<51> ), .clk(clk), .rst(
        n662) );
  dff_60 \reg4[52]  ( .q(\fifo3<52> ), .d(\fifo_next3<52> ), .clk(clk), .rst(
        n661) );
  dff_61 \reg4[53]  ( .q(\fifo3<53> ), .d(\fifo_next3<53> ), .clk(clk), .rst(
        n662) );
  dff_62 \reg4[54]  ( .q(\fifo3<54> ), .d(\fifo_next3<54> ), .clk(clk), .rst(
        n661) );
  dff_63 \reg4[55]  ( .q(\fifo3<55> ), .d(\fifo_next3<55> ), .clk(clk), .rst(
        n662) );
  dff_64 \reg4[56]  ( .q(\fifo3<56> ), .d(\fifo_next3<56> ), .clk(clk), .rst(
        n661) );
  dff_65 \reg4[57]  ( .q(\fifo3<57> ), .d(\fifo_next3<57> ), .clk(clk), .rst(
        n662) );
  dff_66 \reg4[58]  ( .q(\fifo3<58> ), .d(\fifo_next3<58> ), .clk(clk), .rst(
        n661) );
  dff_67 \reg4[59]  ( .q(\fifo3<59> ), .d(\fifo_next3<59> ), .clk(clk), .rst(
        n662) );
  dff_68 \reg4[60]  ( .q(\fifo3<60> ), .d(\fifo_next3<60> ), .clk(clk), .rst(
        n661) );
  dff_69 \reg4[61]  ( .q(\fifo3<61> ), .d(\fifo_next3<61> ), .clk(clk), .rst(
        n662) );
  dff_70 \reg4[62]  ( .q(\fifo3<62> ), .d(\fifo_next3<62> ), .clk(clk), .rst(
        n661) );
  dff_71 \reg4[63]  ( .q(\fifo3<63> ), .d(\fifo_next3<63> ), .clk(clk), .rst(
        n662) );
  fulladder2_1 addr ( .A({\readstate<1> , \readstate<0> }), .B({1'b0, 1'b1}), 
        .SUM({\readstate_plus1<1> , \readstate_plus1<0> }) );
  fulladder2_0 addw ( .A({\writestate<1> , \writestate<0> }), .B({1'b0, 1'b1}), 
        .SUM({\writestate_plus1<1> , \writestate_plus1<0> }) );
  counter5 countrw ( .push(n151), .pop(data_out_valid), .rst(n660), .clk(clk), 
        .currentState({\rwcounter<3> , \rwcounter<2> , \rwcounter<1> , 
        \rwcounter<0> }) );
  dff_6 \rs1[0]  ( .q(\readstate<0> ), .d(\readstate_next<0> ), .clk(clk), 
        .rst(n661) );
  dff_7 \rs1[1]  ( .q(\readstate<1> ), .d(\readstate_next<1> ), .clk(clk), 
        .rst(n662) );
  dff_4 \ws1[0]  ( .q(\writestate<0> ), .d(n664), .clk(clk), .rst(n661) );
  dff_5 \ws1[1]  ( .q(\writestate<1> ), .d(n663), .clk(clk), .rst(n662) );
  INVX2 U219 ( .A(n659), .Y(n660) );
  INVX1 U220 ( .A(\writestate<1> ), .Y(n376) );
  INVX1 U221 ( .A(\fifo0<1> ), .Y(n632) );
  INVX1 U222 ( .A(\fifo0<2> ), .Y(n631) );
  INVX1 U223 ( .A(\fifo0<3> ), .Y(n630) );
  INVX1 U224 ( .A(\fifo0<4> ), .Y(n629) );
  INVX1 U225 ( .A(\fifo0<5> ), .Y(n628) );
  INVX1 U226 ( .A(\fifo0<6> ), .Y(n627) );
  INVX1 U227 ( .A(\fifo0<7> ), .Y(n626) );
  INVX1 U228 ( .A(\fifo0<8> ), .Y(n625) );
  INVX1 U229 ( .A(\fifo0<9> ), .Y(n624) );
  INVX1 U230 ( .A(\fifo0<10> ), .Y(n623) );
  INVX1 U231 ( .A(\fifo0<11> ), .Y(n622) );
  INVX1 U232 ( .A(\fifo0<12> ), .Y(n621) );
  INVX1 U233 ( .A(\fifo0<13> ), .Y(n620) );
  INVX1 U234 ( .A(\fifo0<14> ), .Y(n619) );
  INVX1 U235 ( .A(\fifo0<15> ), .Y(n618) );
  INVX1 U236 ( .A(\fifo0<16> ), .Y(n617) );
  INVX1 U237 ( .A(\fifo0<17> ), .Y(n616) );
  INVX1 U238 ( .A(\fifo0<18> ), .Y(n615) );
  INVX1 U239 ( .A(\fifo0<19> ), .Y(n614) );
  INVX1 U240 ( .A(\fifo0<20> ), .Y(n613) );
  INVX1 U241 ( .A(\fifo0<21> ), .Y(n612) );
  INVX1 U242 ( .A(\fifo0<22> ), .Y(n611) );
  INVX1 U243 ( .A(\fifo0<23> ), .Y(n610) );
  INVX1 U244 ( .A(\fifo0<24> ), .Y(n609) );
  INVX1 U245 ( .A(\fifo0<25> ), .Y(n608) );
  INVX1 U246 ( .A(\fifo0<26> ), .Y(n607) );
  INVX1 U247 ( .A(\fifo0<27> ), .Y(n606) );
  INVX1 U248 ( .A(\fifo0<28> ), .Y(n605) );
  INVX1 U249 ( .A(\fifo0<29> ), .Y(n604) );
  INVX1 U250 ( .A(\fifo0<30> ), .Y(n603) );
  INVX1 U251 ( .A(\fifo0<31> ), .Y(n602) );
  INVX1 U252 ( .A(\fifo0<32> ), .Y(n601) );
  INVX1 U253 ( .A(\fifo0<33> ), .Y(n600) );
  INVX1 U254 ( .A(\fifo0<34> ), .Y(n599) );
  INVX1 U255 ( .A(\fifo0<35> ), .Y(n598) );
  INVX1 U256 ( .A(\fifo0<36> ), .Y(n597) );
  INVX1 U257 ( .A(\fifo0<37> ), .Y(n596) );
  INVX1 U258 ( .A(\fifo0<38> ), .Y(n595) );
  INVX1 U259 ( .A(\fifo0<39> ), .Y(n594) );
  INVX1 U260 ( .A(\fifo0<40> ), .Y(n593) );
  INVX1 U261 ( .A(\fifo0<41> ), .Y(n592) );
  INVX1 U262 ( .A(\fifo0<42> ), .Y(n591) );
  INVX1 U263 ( .A(\fifo0<43> ), .Y(n590) );
  INVX1 U264 ( .A(\fifo0<44> ), .Y(n589) );
  INVX1 U265 ( .A(\fifo0<45> ), .Y(n588) );
  INVX1 U266 ( .A(\fifo0<46> ), .Y(n587) );
  INVX1 U267 ( .A(\fifo0<47> ), .Y(n586) );
  INVX1 U268 ( .A(\fifo0<48> ), .Y(n585) );
  INVX1 U269 ( .A(\fifo0<49> ), .Y(n584) );
  INVX1 U270 ( .A(\fifo0<50> ), .Y(n583) );
  INVX1 U271 ( .A(\fifo0<51> ), .Y(n582) );
  INVX1 U272 ( .A(\fifo0<52> ), .Y(n581) );
  INVX1 U273 ( .A(\fifo0<53> ), .Y(n580) );
  INVX1 U274 ( .A(\fifo0<54> ), .Y(n579) );
  INVX1 U275 ( .A(\fifo0<55> ), .Y(n578) );
  INVX1 U276 ( .A(\fifo0<56> ), .Y(n577) );
  INVX1 U277 ( .A(\fifo0<57> ), .Y(n576) );
  INVX1 U278 ( .A(\fifo0<58> ), .Y(n575) );
  INVX1 U279 ( .A(\fifo0<59> ), .Y(n574) );
  INVX1 U280 ( .A(\fifo0<60> ), .Y(n573) );
  INVX1 U281 ( .A(\fifo0<61> ), .Y(n572) );
  INVX1 U282 ( .A(\fifo0<62> ), .Y(n571) );
  INVX1 U283 ( .A(\fifo0<63> ), .Y(n570) );
  INVX1 U284 ( .A(\fifo1<0> ), .Y(n569) );
  INVX1 U285 ( .A(\fifo1<1> ), .Y(n568) );
  INVX1 U286 ( .A(\fifo1<2> ), .Y(n567) );
  INVX1 U287 ( .A(\fifo1<3> ), .Y(n566) );
  INVX1 U288 ( .A(\fifo1<4> ), .Y(n565) );
  INVX1 U289 ( .A(\fifo1<5> ), .Y(n564) );
  INVX1 U290 ( .A(\fifo1<6> ), .Y(n563) );
  INVX1 U291 ( .A(\fifo1<7> ), .Y(n562) );
  INVX1 U292 ( .A(\fifo1<8> ), .Y(n561) );
  INVX1 U293 ( .A(\fifo1<9> ), .Y(n560) );
  INVX1 U294 ( .A(\fifo1<10> ), .Y(n559) );
  INVX1 U295 ( .A(\fifo1<11> ), .Y(n558) );
  INVX1 U296 ( .A(\fifo1<12> ), .Y(n557) );
  INVX1 U297 ( .A(\fifo1<13> ), .Y(n556) );
  INVX1 U298 ( .A(\fifo1<14> ), .Y(n555) );
  INVX1 U299 ( .A(\fifo1<15> ), .Y(n554) );
  INVX1 U300 ( .A(\fifo1<16> ), .Y(n553) );
  INVX1 U301 ( .A(\fifo1<17> ), .Y(n552) );
  INVX1 U302 ( .A(\fifo1<18> ), .Y(n551) );
  INVX1 U303 ( .A(\fifo1<19> ), .Y(n550) );
  INVX1 U304 ( .A(\fifo1<20> ), .Y(n549) );
  INVX1 U305 ( .A(\fifo1<21> ), .Y(n548) );
  INVX1 U306 ( .A(\fifo1<22> ), .Y(n547) );
  INVX1 U307 ( .A(\fifo1<23> ), .Y(n546) );
  INVX1 U308 ( .A(\fifo1<24> ), .Y(n545) );
  INVX1 U309 ( .A(\fifo1<25> ), .Y(n544) );
  INVX1 U310 ( .A(\fifo1<26> ), .Y(n543) );
  INVX1 U311 ( .A(\fifo1<27> ), .Y(n542) );
  INVX1 U312 ( .A(\fifo1<28> ), .Y(n541) );
  INVX1 U313 ( .A(\fifo1<29> ), .Y(n540) );
  INVX1 U314 ( .A(\fifo1<30> ), .Y(n539) );
  INVX1 U315 ( .A(\fifo1<31> ), .Y(n538) );
  INVX1 U316 ( .A(\fifo1<32> ), .Y(n537) );
  INVX1 U317 ( .A(\fifo1<33> ), .Y(n536) );
  INVX1 U318 ( .A(\fifo1<34> ), .Y(n535) );
  INVX1 U319 ( .A(\fifo1<35> ), .Y(n534) );
  INVX1 U320 ( .A(\fifo1<36> ), .Y(n533) );
  INVX1 U321 ( .A(\fifo1<37> ), .Y(n532) );
  INVX1 U322 ( .A(\fifo1<38> ), .Y(n531) );
  INVX1 U323 ( .A(\fifo1<39> ), .Y(n530) );
  INVX1 U324 ( .A(\fifo1<40> ), .Y(n529) );
  INVX1 U325 ( .A(\fifo1<41> ), .Y(n528) );
  INVX1 U326 ( .A(\fifo1<42> ), .Y(n527) );
  INVX1 U327 ( .A(\fifo1<43> ), .Y(n526) );
  INVX1 U328 ( .A(\fifo1<44> ), .Y(n525) );
  INVX1 U329 ( .A(\fifo1<45> ), .Y(n524) );
  INVX1 U330 ( .A(\fifo1<46> ), .Y(n523) );
  INVX1 U331 ( .A(\fifo1<47> ), .Y(n522) );
  INVX1 U332 ( .A(\fifo1<48> ), .Y(n521) );
  INVX1 U333 ( .A(\fifo1<49> ), .Y(n520) );
  INVX1 U334 ( .A(\fifo1<50> ), .Y(n519) );
  INVX1 U335 ( .A(\fifo1<51> ), .Y(n518) );
  INVX1 U336 ( .A(\fifo1<52> ), .Y(n517) );
  INVX1 U337 ( .A(\fifo1<53> ), .Y(n516) );
  INVX1 U338 ( .A(\fifo1<54> ), .Y(n515) );
  INVX1 U339 ( .A(\fifo1<55> ), .Y(n514) );
  INVX1 U340 ( .A(\fifo1<56> ), .Y(n513) );
  INVX1 U341 ( .A(\fifo1<57> ), .Y(n512) );
  INVX1 U342 ( .A(\fifo1<58> ), .Y(n511) );
  INVX1 U343 ( .A(\fifo1<59> ), .Y(n510) );
  INVX1 U344 ( .A(\fifo1<60> ), .Y(n509) );
  INVX1 U345 ( .A(\fifo1<61> ), .Y(n508) );
  INVX1 U346 ( .A(\fifo1<62> ), .Y(n507) );
  INVX1 U347 ( .A(\fifo1<63> ), .Y(n506) );
  INVX1 U348 ( .A(\fifo2<0> ), .Y(n505) );
  INVX1 U349 ( .A(\fifo2<1> ), .Y(n504) );
  INVX1 U350 ( .A(\fifo2<2> ), .Y(n503) );
  INVX1 U351 ( .A(\fifo2<3> ), .Y(n502) );
  INVX1 U352 ( .A(\fifo2<4> ), .Y(n501) );
  INVX1 U353 ( .A(\fifo2<5> ), .Y(n500) );
  INVX1 U354 ( .A(\fifo2<6> ), .Y(n499) );
  INVX1 U355 ( .A(\fifo2<7> ), .Y(n498) );
  INVX1 U356 ( .A(\fifo2<8> ), .Y(n497) );
  INVX1 U357 ( .A(\fifo2<9> ), .Y(n496) );
  INVX1 U358 ( .A(\fifo2<10> ), .Y(n495) );
  INVX1 U359 ( .A(\fifo2<11> ), .Y(n494) );
  INVX1 U360 ( .A(\fifo2<12> ), .Y(n493) );
  INVX1 U361 ( .A(\fifo2<13> ), .Y(n492) );
  INVX1 U362 ( .A(\fifo2<14> ), .Y(n491) );
  INVX1 U363 ( .A(\fifo2<15> ), .Y(n490) );
  INVX1 U364 ( .A(\fifo2<16> ), .Y(n489) );
  INVX1 U365 ( .A(\fifo2<17> ), .Y(n488) );
  INVX1 U366 ( .A(\fifo2<18> ), .Y(n487) );
  INVX1 U367 ( .A(\fifo2<19> ), .Y(n486) );
  INVX1 U368 ( .A(\fifo2<20> ), .Y(n485) );
  INVX1 U369 ( .A(\fifo2<21> ), .Y(n484) );
  INVX1 U370 ( .A(\fifo2<22> ), .Y(n483) );
  INVX1 U371 ( .A(\fifo2<23> ), .Y(n482) );
  INVX1 U372 ( .A(\fifo2<24> ), .Y(n481) );
  INVX1 U373 ( .A(\fifo2<25> ), .Y(n480) );
  INVX1 U374 ( .A(\fifo2<26> ), .Y(n479) );
  INVX1 U375 ( .A(\fifo2<27> ), .Y(n478) );
  INVX1 U376 ( .A(\fifo2<28> ), .Y(n477) );
  INVX1 U377 ( .A(\fifo2<29> ), .Y(n476) );
  INVX1 U378 ( .A(\fifo2<30> ), .Y(n475) );
  INVX1 U379 ( .A(\fifo2<31> ), .Y(n474) );
  INVX1 U380 ( .A(\fifo2<32> ), .Y(n473) );
  INVX1 U381 ( .A(\fifo2<33> ), .Y(n472) );
  INVX1 U382 ( .A(\fifo2<34> ), .Y(n471) );
  INVX1 U383 ( .A(\fifo2<35> ), .Y(n470) );
  INVX1 U384 ( .A(\fifo2<36> ), .Y(n469) );
  INVX1 U385 ( .A(\fifo2<37> ), .Y(n468) );
  INVX1 U386 ( .A(\fifo2<38> ), .Y(n467) );
  INVX1 U387 ( .A(\fifo2<39> ), .Y(n466) );
  INVX1 U388 ( .A(\fifo2<40> ), .Y(n465) );
  INVX1 U389 ( .A(\fifo2<41> ), .Y(n464) );
  INVX1 U390 ( .A(\fifo2<42> ), .Y(n463) );
  INVX1 U391 ( .A(\fifo2<43> ), .Y(n462) );
  INVX1 U392 ( .A(\fifo2<44> ), .Y(n461) );
  INVX1 U393 ( .A(\fifo2<45> ), .Y(n460) );
  INVX1 U394 ( .A(\fifo2<46> ), .Y(n459) );
  INVX1 U395 ( .A(\fifo2<47> ), .Y(n458) );
  INVX1 U396 ( .A(\fifo2<48> ), .Y(n457) );
  INVX1 U397 ( .A(\fifo2<49> ), .Y(n456) );
  INVX1 U398 ( .A(\fifo2<50> ), .Y(n455) );
  INVX1 U399 ( .A(\fifo2<51> ), .Y(n454) );
  INVX1 U400 ( .A(\fifo2<52> ), .Y(n453) );
  INVX1 U401 ( .A(\fifo2<53> ), .Y(n452) );
  INVX1 U402 ( .A(\fifo2<54> ), .Y(n451) );
  INVX1 U403 ( .A(\fifo2<55> ), .Y(n450) );
  INVX1 U404 ( .A(\fifo2<56> ), .Y(n449) );
  INVX1 U405 ( .A(\fifo2<57> ), .Y(n448) );
  INVX1 U406 ( .A(\fifo2<58> ), .Y(n447) );
  INVX1 U407 ( .A(\fifo2<59> ), .Y(n446) );
  INVX1 U408 ( .A(\fifo2<60> ), .Y(n445) );
  INVX1 U409 ( .A(\fifo2<61> ), .Y(n444) );
  INVX1 U410 ( .A(\fifo2<62> ), .Y(n443) );
  INVX1 U411 ( .A(\fifo2<63> ), .Y(n442) );
  INVX1 U412 ( .A(\fifo3<0> ), .Y(n441) );
  INVX1 U413 ( .A(\data_in<1> ), .Y(n312) );
  INVX1 U414 ( .A(\fifo3<1> ), .Y(n440) );
  INVX1 U415 ( .A(\data_in<2> ), .Y(n313) );
  INVX1 U416 ( .A(\fifo3<2> ), .Y(n439) );
  INVX1 U417 ( .A(\data_in<3> ), .Y(n314) );
  INVX1 U418 ( .A(\fifo3<3> ), .Y(n438) );
  INVX1 U419 ( .A(\data_in<4> ), .Y(n315) );
  INVX1 U420 ( .A(\fifo3<4> ), .Y(n437) );
  INVX1 U421 ( .A(\data_in<5> ), .Y(n316) );
  INVX1 U422 ( .A(\fifo3<5> ), .Y(n436) );
  INVX1 U423 ( .A(\data_in<6> ), .Y(n317) );
  INVX1 U424 ( .A(\fifo3<6> ), .Y(n435) );
  INVX1 U425 ( .A(\data_in<7> ), .Y(n318) );
  INVX1 U426 ( .A(\fifo3<7> ), .Y(n434) );
  INVX1 U427 ( .A(\data_in<8> ), .Y(n319) );
  INVX1 U428 ( .A(\fifo3<8> ), .Y(n433) );
  INVX1 U429 ( .A(\data_in<9> ), .Y(n320) );
  INVX1 U430 ( .A(\fifo3<9> ), .Y(n432) );
  INVX1 U431 ( .A(\data_in<10> ), .Y(n321) );
  INVX1 U432 ( .A(\fifo3<10> ), .Y(n431) );
  INVX1 U433 ( .A(\data_in<11> ), .Y(n322) );
  INVX1 U434 ( .A(\fifo3<11> ), .Y(n430) );
  INVX1 U435 ( .A(\data_in<12> ), .Y(n323) );
  INVX1 U436 ( .A(\fifo3<12> ), .Y(n429) );
  INVX1 U437 ( .A(\data_in<13> ), .Y(n324) );
  INVX1 U438 ( .A(\fifo3<13> ), .Y(n428) );
  INVX1 U439 ( .A(\data_in<14> ), .Y(n325) );
  INVX1 U440 ( .A(\fifo3<14> ), .Y(n427) );
  INVX1 U441 ( .A(\data_in<15> ), .Y(n326) );
  INVX1 U442 ( .A(\fifo3<15> ), .Y(n426) );
  INVX1 U443 ( .A(\data_in<16> ), .Y(n327) );
  INVX1 U444 ( .A(\fifo3<16> ), .Y(n425) );
  INVX1 U445 ( .A(\data_in<17> ), .Y(n328) );
  INVX1 U446 ( .A(\fifo3<17> ), .Y(n424) );
  INVX1 U447 ( .A(\data_in<18> ), .Y(n329) );
  INVX1 U448 ( .A(\fifo3<18> ), .Y(n423) );
  INVX1 U449 ( .A(\data_in<19> ), .Y(n330) );
  INVX1 U450 ( .A(\fifo3<19> ), .Y(n422) );
  INVX1 U451 ( .A(\data_in<20> ), .Y(n331) );
  INVX1 U452 ( .A(\fifo3<20> ), .Y(n421) );
  INVX1 U453 ( .A(\data_in<21> ), .Y(n332) );
  INVX1 U454 ( .A(\fifo3<21> ), .Y(n420) );
  INVX1 U455 ( .A(\data_in<22> ), .Y(n333) );
  INVX1 U456 ( .A(\fifo3<22> ), .Y(n419) );
  INVX1 U457 ( .A(\data_in<23> ), .Y(n334) );
  INVX1 U458 ( .A(\fifo3<23> ), .Y(n418) );
  INVX1 U459 ( .A(\data_in<24> ), .Y(n335) );
  INVX1 U460 ( .A(\fifo3<24> ), .Y(n417) );
  INVX1 U461 ( .A(\data_in<25> ), .Y(n336) );
  INVX1 U462 ( .A(\fifo3<25> ), .Y(n416) );
  INVX1 U463 ( .A(\data_in<26> ), .Y(n337) );
  INVX1 U464 ( .A(\fifo3<26> ), .Y(n415) );
  INVX1 U465 ( .A(\data_in<27> ), .Y(n338) );
  INVX1 U466 ( .A(\fifo3<27> ), .Y(n414) );
  INVX1 U467 ( .A(\data_in<28> ), .Y(n339) );
  INVX1 U468 ( .A(\fifo3<28> ), .Y(n413) );
  INVX1 U469 ( .A(\data_in<29> ), .Y(n340) );
  INVX1 U470 ( .A(\fifo3<29> ), .Y(n412) );
  INVX1 U471 ( .A(\data_in<30> ), .Y(n341) );
  INVX1 U472 ( .A(\fifo3<30> ), .Y(n411) );
  INVX1 U473 ( .A(\data_in<31> ), .Y(n342) );
  INVX1 U474 ( .A(\fifo3<31> ), .Y(n410) );
  INVX1 U475 ( .A(\data_in<32> ), .Y(n343) );
  INVX1 U476 ( .A(\fifo3<32> ), .Y(n409) );
  INVX1 U477 ( .A(\data_in<33> ), .Y(n344) );
  INVX1 U478 ( .A(\fifo3<33> ), .Y(n408) );
  INVX1 U479 ( .A(\data_in<34> ), .Y(n345) );
  INVX1 U480 ( .A(\fifo3<34> ), .Y(n407) );
  INVX1 U481 ( .A(\data_in<35> ), .Y(n346) );
  INVX1 U482 ( .A(\fifo3<35> ), .Y(n406) );
  INVX1 U483 ( .A(\data_in<36> ), .Y(n347) );
  INVX1 U484 ( .A(\fifo3<36> ), .Y(n405) );
  INVX1 U485 ( .A(\data_in<37> ), .Y(n348) );
  INVX1 U486 ( .A(\fifo3<37> ), .Y(n404) );
  INVX1 U487 ( .A(\data_in<38> ), .Y(n349) );
  INVX1 U488 ( .A(\fifo3<38> ), .Y(n403) );
  INVX1 U489 ( .A(\data_in<39> ), .Y(n350) );
  INVX1 U490 ( .A(\fifo3<39> ), .Y(n402) );
  INVX1 U491 ( .A(\data_in<40> ), .Y(n351) );
  INVX1 U492 ( .A(\fifo3<40> ), .Y(n401) );
  INVX1 U493 ( .A(\data_in<41> ), .Y(n352) );
  INVX1 U494 ( .A(\fifo3<41> ), .Y(n400) );
  INVX1 U495 ( .A(\data_in<42> ), .Y(n353) );
  INVX1 U496 ( .A(\fifo3<42> ), .Y(n399) );
  INVX1 U497 ( .A(\data_in<43> ), .Y(n354) );
  INVX1 U498 ( .A(\fifo3<43> ), .Y(n398) );
  INVX1 U499 ( .A(\data_in<44> ), .Y(n355) );
  INVX1 U500 ( .A(\fifo3<44> ), .Y(n397) );
  INVX1 U501 ( .A(\data_in<45> ), .Y(n356) );
  INVX1 U502 ( .A(\fifo3<45> ), .Y(n396) );
  INVX1 U503 ( .A(\data_in<46> ), .Y(n357) );
  INVX1 U504 ( .A(\fifo3<46> ), .Y(n395) );
  INVX1 U505 ( .A(\data_in<47> ), .Y(n358) );
  INVX1 U506 ( .A(\fifo3<47> ), .Y(n394) );
  INVX1 U507 ( .A(\data_in<48> ), .Y(n359) );
  INVX1 U508 ( .A(\fifo3<48> ), .Y(n393) );
  INVX1 U509 ( .A(\data_in<49> ), .Y(n360) );
  INVX1 U510 ( .A(\fifo3<49> ), .Y(n392) );
  INVX1 U511 ( .A(\data_in<50> ), .Y(n361) );
  INVX1 U512 ( .A(\fifo3<50> ), .Y(n391) );
  INVX1 U513 ( .A(\data_in<51> ), .Y(n362) );
  INVX1 U514 ( .A(\fifo3<51> ), .Y(n390) );
  INVX1 U515 ( .A(\data_in<52> ), .Y(n363) );
  INVX1 U516 ( .A(\fifo3<52> ), .Y(n389) );
  INVX1 U517 ( .A(\data_in<53> ), .Y(n364) );
  INVX1 U518 ( .A(\fifo3<53> ), .Y(n388) );
  INVX1 U519 ( .A(\data_in<54> ), .Y(n365) );
  INVX1 U520 ( .A(\fifo3<54> ), .Y(n387) );
  INVX1 U521 ( .A(\data_in<55> ), .Y(n366) );
  INVX1 U522 ( .A(\fifo3<55> ), .Y(n386) );
  INVX1 U523 ( .A(\data_in<56> ), .Y(n367) );
  INVX1 U524 ( .A(\fifo3<56> ), .Y(n385) );
  INVX1 U525 ( .A(\data_in<57> ), .Y(n368) );
  INVX1 U526 ( .A(\fifo3<57> ), .Y(n384) );
  INVX1 U527 ( .A(\data_in<58> ), .Y(n369) );
  INVX1 U528 ( .A(\fifo3<58> ), .Y(n383) );
  INVX1 U529 ( .A(\data_in<59> ), .Y(n370) );
  INVX1 U530 ( .A(\fifo3<59> ), .Y(n382) );
  INVX1 U531 ( .A(\data_in<60> ), .Y(n371) );
  INVX1 U532 ( .A(\fifo3<60> ), .Y(n381) );
  INVX1 U533 ( .A(\data_in<61> ), .Y(n372) );
  INVX1 U534 ( .A(\fifo3<61> ), .Y(n380) );
  INVX1 U535 ( .A(\data_in<62> ), .Y(n373) );
  INVX1 U536 ( .A(\fifo3<62> ), .Y(n379) );
  INVX1 U537 ( .A(\data_in<63> ), .Y(n374) );
  INVX1 U538 ( .A(\fifo3<63> ), .Y(n378) );
  INVX1 U539 ( .A(\readstate<0> ), .Y(n665) );
  INVX1 U540 ( .A(\readstate<1> ), .Y(n666) );
  INVX1 U541 ( .A(\data_in<0> ), .Y(n311) );
  INVX1 U542 ( .A(\fifo0<0> ), .Y(n375) );
  AND2X1 U543 ( .A(pop_fifo), .B(n299), .Y(data_out_valid) );
  AND2X1 U544 ( .A(data_in_valid), .B(n303), .Y(n151) );
  INVX1 U545 ( .A(\writestate<0> ), .Y(n377) );
  AND2X1 U546 ( .A(\writestate<1> ), .B(n306), .Y(n301) );
  AND2X1 U547 ( .A(n306), .B(n376), .Y(n304) );
  INVX1 U548 ( .A(\rwcounter<2> ), .Y(n667) );
  INVX1 U549 ( .A(n289), .Y(n638) );
  INVX1 U550 ( .A(n289), .Y(n637) );
  INVX1 U551 ( .A(n288), .Y(n643) );
  INVX1 U552 ( .A(n288), .Y(n644) );
  INVX1 U553 ( .A(n290), .Y(n641) );
  INVX1 U554 ( .A(n290), .Y(n640) );
  INVX1 U555 ( .A(n287), .Y(n635) );
  INVX1 U556 ( .A(n287), .Y(n634) );
  INVX2 U557 ( .A(n659), .Y(n661) );
  INVX2 U558 ( .A(n659), .Y(n662) );
  INVX1 U559 ( .A(n647), .Y(n645) );
  AND2X1 U560 ( .A(n665), .B(n666), .Y(n23) );
  INVX1 U561 ( .A(n23), .Y(n647) );
  AND2X1 U562 ( .A(\rwcounter<2> ), .B(n16), .Y(fifo_full) );
  AND2X1 U563 ( .A(n16), .B(n667), .Y(fifo_empty) );
  INVX1 U564 ( .A(n21), .Y(n655) );
  AND2X1 U565 ( .A(\readstate<0> ), .B(\readstate<1> ), .Y(n20) );
  INVX1 U566 ( .A(n20), .Y(n658) );
  AND2X1 U567 ( .A(\readstate<0> ), .B(n666), .Y(n22) );
  INVX1 U568 ( .A(n22), .Y(n651) );
  INVX1 U569 ( .A(n287), .Y(n633) );
  INVX1 U570 ( .A(n288), .Y(n642) );
  INVX1 U571 ( .A(n290), .Y(n639) );
  INVX1 U572 ( .A(n289), .Y(n636) );
  INVX1 U573 ( .A(n647), .Y(n646) );
  AND2X1 U574 ( .A(\readstate<1> ), .B(n665), .Y(n21) );
  INVX1 U575 ( .A(rst), .Y(n659) );
  INVX1 U576 ( .A(n151), .Y(n152) );
  INVX1 U577 ( .A(n655), .Y(n654) );
  INVX1 U578 ( .A(n651), .Y(n650) );
  INVX1 U579 ( .A(n655), .Y(n653) );
  INVX1 U580 ( .A(n658), .Y(n657) );
  INVX1 U581 ( .A(n651), .Y(n649) );
  INVX1 U582 ( .A(n655), .Y(n652) );
  INVX1 U583 ( .A(n651), .Y(n648) );
  INVX1 U584 ( .A(n658), .Y(n656) );
  AND2X1 U585 ( .A(\readstate_plus1<0> ), .B(data_out_valid), .Y(n153) );
  INVX1 U586 ( .A(n153), .Y(n154) );
  AND2X1 U587 ( .A(\readstate_plus1<1> ), .B(data_out_valid), .Y(n155) );
  INVX1 U588 ( .A(n155), .Y(n156) );
  BUFX2 U589 ( .A(n149), .Y(n157) );
  BUFX2 U590 ( .A(n147), .Y(n158) );
  BUFX2 U591 ( .A(n145), .Y(n159) );
  BUFX2 U592 ( .A(n143), .Y(n160) );
  BUFX2 U593 ( .A(n141), .Y(n161) );
  BUFX2 U594 ( .A(n139), .Y(n162) );
  BUFX2 U595 ( .A(n137), .Y(n163) );
  BUFX2 U596 ( .A(n135), .Y(n164) );
  BUFX2 U597 ( .A(n133), .Y(n165) );
  BUFX2 U598 ( .A(n131), .Y(n166) );
  BUFX2 U599 ( .A(n129), .Y(n167) );
  BUFX2 U600 ( .A(n127), .Y(n168) );
  BUFX2 U601 ( .A(n125), .Y(n169) );
  BUFX2 U602 ( .A(n123), .Y(n170) );
  BUFX2 U603 ( .A(n121), .Y(n171) );
  BUFX2 U604 ( .A(n119), .Y(n172) );
  BUFX2 U605 ( .A(n117), .Y(n173) );
  BUFX2 U606 ( .A(n115), .Y(n174) );
  BUFX2 U607 ( .A(n113), .Y(n175) );
  BUFX2 U608 ( .A(n111), .Y(n176) );
  BUFX2 U609 ( .A(n109), .Y(n177) );
  BUFX2 U610 ( .A(n107), .Y(n178) );
  BUFX2 U611 ( .A(n105), .Y(n179) );
  BUFX2 U612 ( .A(n103), .Y(n180) );
  BUFX2 U613 ( .A(n101), .Y(n181) );
  BUFX2 U614 ( .A(n99), .Y(n182) );
  BUFX2 U615 ( .A(n97), .Y(n183) );
  BUFX2 U616 ( .A(n95), .Y(n184) );
  BUFX2 U617 ( .A(n93), .Y(n185) );
  BUFX2 U618 ( .A(n91), .Y(n186) );
  BUFX2 U619 ( .A(n89), .Y(n187) );
  BUFX2 U620 ( .A(n87), .Y(n188) );
  BUFX2 U621 ( .A(n85), .Y(n189) );
  BUFX2 U622 ( .A(n83), .Y(n190) );
  BUFX2 U623 ( .A(n81), .Y(n191) );
  BUFX2 U624 ( .A(n79), .Y(n192) );
  BUFX2 U625 ( .A(n77), .Y(n193) );
  BUFX2 U626 ( .A(n75), .Y(n194) );
  BUFX2 U627 ( .A(n73), .Y(n195) );
  BUFX2 U628 ( .A(n71), .Y(n196) );
  BUFX2 U629 ( .A(n69), .Y(n197) );
  BUFX2 U630 ( .A(n67), .Y(n198) );
  BUFX2 U631 ( .A(n65), .Y(n199) );
  BUFX2 U632 ( .A(n63), .Y(n200) );
  BUFX2 U633 ( .A(n61), .Y(n201) );
  BUFX2 U634 ( .A(n59), .Y(n202) );
  BUFX2 U635 ( .A(n57), .Y(n203) );
  BUFX2 U636 ( .A(n55), .Y(n204) );
  BUFX2 U637 ( .A(n53), .Y(n205) );
  BUFX2 U638 ( .A(n51), .Y(n206) );
  BUFX2 U639 ( .A(n49), .Y(n207) );
  BUFX2 U640 ( .A(n47), .Y(n208) );
  BUFX2 U641 ( .A(n45), .Y(n209) );
  BUFX2 U642 ( .A(n43), .Y(n210) );
  BUFX2 U643 ( .A(n41), .Y(n211) );
  BUFX2 U644 ( .A(n39), .Y(n212) );
  BUFX2 U645 ( .A(n37), .Y(n213) );
  BUFX2 U646 ( .A(n35), .Y(n214) );
  BUFX2 U647 ( .A(n33), .Y(n215) );
  BUFX2 U648 ( .A(n31), .Y(n216) );
  BUFX2 U649 ( .A(n29), .Y(n217) );
  BUFX2 U650 ( .A(n27), .Y(n218) );
  BUFX2 U651 ( .A(n25), .Y(n219) );
  BUFX2 U652 ( .A(n19), .Y(n220) );
  BUFX2 U653 ( .A(n148), .Y(n221) );
  BUFX2 U654 ( .A(n146), .Y(n222) );
  BUFX2 U655 ( .A(n144), .Y(n223) );
  BUFX2 U656 ( .A(n142), .Y(n224) );
  BUFX2 U657 ( .A(n140), .Y(n225) );
  BUFX2 U658 ( .A(n138), .Y(n226) );
  BUFX2 U659 ( .A(n136), .Y(n227) );
  BUFX2 U660 ( .A(n134), .Y(n228) );
  BUFX2 U661 ( .A(n132), .Y(n229) );
  BUFX2 U662 ( .A(n130), .Y(n230) );
  BUFX2 U663 ( .A(n128), .Y(n231) );
  BUFX2 U664 ( .A(n126), .Y(n232) );
  BUFX2 U665 ( .A(n124), .Y(n233) );
  BUFX2 U666 ( .A(n122), .Y(n234) );
  BUFX2 U667 ( .A(n120), .Y(n235) );
  BUFX2 U668 ( .A(n118), .Y(n236) );
  BUFX2 U669 ( .A(n116), .Y(n237) );
  BUFX2 U670 ( .A(n114), .Y(n238) );
  BUFX2 U671 ( .A(n112), .Y(n239) );
  BUFX2 U672 ( .A(n110), .Y(n240) );
  BUFX2 U673 ( .A(n108), .Y(n241) );
  BUFX2 U674 ( .A(n106), .Y(n242) );
  BUFX2 U675 ( .A(n104), .Y(n243) );
  BUFX2 U676 ( .A(n102), .Y(n244) );
  BUFX2 U677 ( .A(n100), .Y(n245) );
  BUFX2 U678 ( .A(n98), .Y(n246) );
  BUFX2 U679 ( .A(n96), .Y(n247) );
  BUFX2 U680 ( .A(n94), .Y(n248) );
  BUFX2 U681 ( .A(n92), .Y(n249) );
  BUFX2 U682 ( .A(n90), .Y(n250) );
  BUFX2 U683 ( .A(n88), .Y(n251) );
  BUFX2 U684 ( .A(n86), .Y(n252) );
  BUFX2 U685 ( .A(n84), .Y(n253) );
  BUFX2 U686 ( .A(n82), .Y(n254) );
  BUFX2 U687 ( .A(n80), .Y(n255) );
  BUFX2 U688 ( .A(n78), .Y(n256) );
  BUFX2 U689 ( .A(n76), .Y(n257) );
  BUFX2 U690 ( .A(n74), .Y(n258) );
  BUFX2 U691 ( .A(n72), .Y(n259) );
  BUFX2 U692 ( .A(n70), .Y(n260) );
  BUFX2 U693 ( .A(n68), .Y(n261) );
  BUFX2 U694 ( .A(n66), .Y(n262) );
  BUFX2 U695 ( .A(n64), .Y(n263) );
  BUFX2 U696 ( .A(n62), .Y(n264) );
  BUFX2 U697 ( .A(n60), .Y(n265) );
  BUFX2 U698 ( .A(n58), .Y(n266) );
  BUFX2 U699 ( .A(n56), .Y(n267) );
  BUFX2 U700 ( .A(n54), .Y(n268) );
  BUFX2 U701 ( .A(n52), .Y(n269) );
  BUFX2 U702 ( .A(n50), .Y(n270) );
  BUFX2 U703 ( .A(n48), .Y(n271) );
  BUFX2 U704 ( .A(n46), .Y(n272) );
  BUFX2 U705 ( .A(n44), .Y(n273) );
  BUFX2 U706 ( .A(n42), .Y(n274) );
  BUFX2 U707 ( .A(n40), .Y(n275) );
  BUFX2 U708 ( .A(n38), .Y(n276) );
  BUFX2 U709 ( .A(n36), .Y(n277) );
  BUFX2 U710 ( .A(n34), .Y(n278) );
  BUFX2 U711 ( .A(n32), .Y(n279) );
  BUFX2 U712 ( .A(n30), .Y(n280) );
  BUFX2 U713 ( .A(n28), .Y(n281) );
  BUFX2 U714 ( .A(n26), .Y(n282) );
  BUFX2 U715 ( .A(n24), .Y(n283) );
  BUFX2 U716 ( .A(n18), .Y(n284) );
  BUFX2 U717 ( .A(n12), .Y(n285) );
  INVX1 U718 ( .A(n285), .Y(n664) );
  BUFX2 U719 ( .A(n10), .Y(n286) );
  INVX1 U720 ( .A(n286), .Y(n663) );
  BUFX2 U721 ( .A(n307), .Y(n287) );
  BUFX2 U722 ( .A(n308), .Y(n288) );
  BUFX2 U723 ( .A(n309), .Y(n289) );
  BUFX2 U724 ( .A(n310), .Y(n290) );
  OR2X1 U725 ( .A(n302), .B(n377), .Y(n291) );
  INVX1 U726 ( .A(n291), .Y(n292) );
  OR2X1 U727 ( .A(\writestate<0> ), .B(n302), .Y(n293) );
  INVX1 U728 ( .A(n293), .Y(n294) );
  OR2X1 U729 ( .A(n377), .B(n305), .Y(n295) );
  INVX1 U730 ( .A(n295), .Y(n296) );
  OR2X1 U731 ( .A(\writestate<0> ), .B(n305), .Y(n297) );
  INVX1 U732 ( .A(n297), .Y(n298) );
  INVX1 U733 ( .A(fifo_empty), .Y(n299) );
  INVX1 U734 ( .A(n301), .Y(n302) );
  INVX1 U735 ( .A(fifo_full), .Y(n303) );
  INVX1 U736 ( .A(n304), .Y(n305) );
  INVX1 U737 ( .A(n152), .Y(n306) );
  MUX2X1 U738 ( .B(n441), .A(n311), .S(n292), .Y(\fifo_next3<0> ) );
  MUX2X1 U739 ( .B(n440), .A(n312), .S(n635), .Y(\fifo_next3<1> ) );
  MUX2X1 U740 ( .B(n439), .A(n313), .S(n635), .Y(\fifo_next3<2> ) );
  MUX2X1 U741 ( .B(n438), .A(n314), .S(n635), .Y(\fifo_next3<3> ) );
  MUX2X1 U742 ( .B(n437), .A(n315), .S(n635), .Y(\fifo_next3<4> ) );
  MUX2X1 U743 ( .B(n436), .A(n316), .S(n635), .Y(\fifo_next3<5> ) );
  MUX2X1 U744 ( .B(n435), .A(n317), .S(n635), .Y(\fifo_next3<6> ) );
  MUX2X1 U745 ( .B(n434), .A(n318), .S(n635), .Y(\fifo_next3<7> ) );
  MUX2X1 U746 ( .B(n433), .A(n319), .S(n635), .Y(\fifo_next3<8> ) );
  MUX2X1 U747 ( .B(n432), .A(n320), .S(n635), .Y(\fifo_next3<9> ) );
  MUX2X1 U748 ( .B(n431), .A(n321), .S(n635), .Y(\fifo_next3<10> ) );
  MUX2X1 U749 ( .B(n430), .A(n322), .S(n635), .Y(\fifo_next3<11> ) );
  MUX2X1 U750 ( .B(n429), .A(n323), .S(n635), .Y(\fifo_next3<12> ) );
  MUX2X1 U751 ( .B(n428), .A(n324), .S(n634), .Y(\fifo_next3<13> ) );
  MUX2X1 U752 ( .B(n427), .A(n325), .S(n634), .Y(\fifo_next3<14> ) );
  MUX2X1 U753 ( .B(n426), .A(n326), .S(n634), .Y(\fifo_next3<15> ) );
  MUX2X1 U754 ( .B(n425), .A(n327), .S(n634), .Y(\fifo_next3<16> ) );
  MUX2X1 U755 ( .B(n424), .A(n328), .S(n634), .Y(\fifo_next3<17> ) );
  MUX2X1 U756 ( .B(n423), .A(n329), .S(n634), .Y(\fifo_next3<18> ) );
  MUX2X1 U757 ( .B(n422), .A(n330), .S(n634), .Y(\fifo_next3<19> ) );
  MUX2X1 U758 ( .B(n421), .A(n331), .S(n634), .Y(\fifo_next3<20> ) );
  MUX2X1 U759 ( .B(n420), .A(n332), .S(n634), .Y(\fifo_next3<21> ) );
  MUX2X1 U760 ( .B(n419), .A(n333), .S(n634), .Y(\fifo_next3<22> ) );
  MUX2X1 U761 ( .B(n418), .A(n334), .S(n634), .Y(\fifo_next3<23> ) );
  MUX2X1 U762 ( .B(n417), .A(n335), .S(n634), .Y(\fifo_next3<24> ) );
  MUX2X1 U763 ( .B(n416), .A(n336), .S(n634), .Y(\fifo_next3<25> ) );
  MUX2X1 U764 ( .B(n415), .A(n337), .S(n635), .Y(\fifo_next3<26> ) );
  MUX2X1 U765 ( .B(n414), .A(n338), .S(n634), .Y(\fifo_next3<27> ) );
  MUX2X1 U766 ( .B(n413), .A(n339), .S(n635), .Y(\fifo_next3<28> ) );
  MUX2X1 U767 ( .B(n412), .A(n340), .S(n634), .Y(\fifo_next3<29> ) );
  MUX2X1 U768 ( .B(n411), .A(n341), .S(n635), .Y(\fifo_next3<30> ) );
  MUX2X1 U769 ( .B(n410), .A(n342), .S(n634), .Y(\fifo_next3<31> ) );
  MUX2X1 U770 ( .B(n409), .A(n343), .S(n635), .Y(\fifo_next3<32> ) );
  MUX2X1 U771 ( .B(n408), .A(n344), .S(n634), .Y(\fifo_next3<33> ) );
  MUX2X1 U772 ( .B(n407), .A(n345), .S(n635), .Y(\fifo_next3<34> ) );
  MUX2X1 U773 ( .B(n406), .A(n346), .S(n634), .Y(\fifo_next3<35> ) );
  MUX2X1 U774 ( .B(n405), .A(n347), .S(n635), .Y(\fifo_next3<36> ) );
  MUX2X1 U775 ( .B(n404), .A(n348), .S(n634), .Y(\fifo_next3<37> ) );
  MUX2X1 U776 ( .B(n403), .A(n349), .S(n633), .Y(\fifo_next3<38> ) );
  MUX2X1 U777 ( .B(n402), .A(n350), .S(n635), .Y(\fifo_next3<39> ) );
  MUX2X1 U778 ( .B(n401), .A(n351), .S(n634), .Y(\fifo_next3<40> ) );
  MUX2X1 U779 ( .B(n400), .A(n352), .S(n633), .Y(\fifo_next3<41> ) );
  MUX2X1 U780 ( .B(n399), .A(n353), .S(n635), .Y(\fifo_next3<42> ) );
  MUX2X1 U781 ( .B(n398), .A(n354), .S(n634), .Y(\fifo_next3<43> ) );
  MUX2X1 U782 ( .B(n397), .A(n355), .S(n633), .Y(\fifo_next3<44> ) );
  MUX2X1 U783 ( .B(n396), .A(n356), .S(n633), .Y(\fifo_next3<45> ) );
  MUX2X1 U784 ( .B(n395), .A(n357), .S(n633), .Y(\fifo_next3<46> ) );
  MUX2X1 U785 ( .B(n394), .A(n358), .S(n633), .Y(\fifo_next3<47> ) );
  MUX2X1 U786 ( .B(n393), .A(n359), .S(n633), .Y(\fifo_next3<48> ) );
  MUX2X1 U787 ( .B(n392), .A(n360), .S(n633), .Y(\fifo_next3<49> ) );
  MUX2X1 U788 ( .B(n391), .A(n361), .S(n633), .Y(\fifo_next3<50> ) );
  MUX2X1 U789 ( .B(n390), .A(n362), .S(n633), .Y(\fifo_next3<51> ) );
  MUX2X1 U790 ( .B(n389), .A(n363), .S(n633), .Y(\fifo_next3<52> ) );
  MUX2X1 U791 ( .B(n388), .A(n364), .S(n633), .Y(\fifo_next3<53> ) );
  MUX2X1 U792 ( .B(n387), .A(n365), .S(n633), .Y(\fifo_next3<54> ) );
  MUX2X1 U793 ( .B(n386), .A(n366), .S(n633), .Y(\fifo_next3<55> ) );
  MUX2X1 U794 ( .B(n385), .A(n367), .S(n633), .Y(\fifo_next3<56> ) );
  MUX2X1 U795 ( .B(n384), .A(n368), .S(n633), .Y(\fifo_next3<57> ) );
  MUX2X1 U796 ( .B(n383), .A(n369), .S(n633), .Y(\fifo_next3<58> ) );
  MUX2X1 U797 ( .B(n382), .A(n370), .S(n633), .Y(\fifo_next3<59> ) );
  MUX2X1 U798 ( .B(n381), .A(n371), .S(n633), .Y(\fifo_next3<60> ) );
  MUX2X1 U799 ( .B(n380), .A(n372), .S(n633), .Y(\fifo_next3<61> ) );
  MUX2X1 U800 ( .B(n379), .A(n373), .S(n633), .Y(\fifo_next3<62> ) );
  MUX2X1 U801 ( .B(n378), .A(n374), .S(n633), .Y(\fifo_next3<63> ) );
  MUX2X1 U802 ( .B(n505), .A(n311), .S(n294), .Y(\fifo_next2<0> ) );
  MUX2X1 U803 ( .B(n504), .A(n312), .S(n644), .Y(\fifo_next2<1> ) );
  MUX2X1 U804 ( .B(n503), .A(n313), .S(n644), .Y(\fifo_next2<2> ) );
  MUX2X1 U805 ( .B(n502), .A(n314), .S(n644), .Y(\fifo_next2<3> ) );
  MUX2X1 U806 ( .B(n501), .A(n315), .S(n644), .Y(\fifo_next2<4> ) );
  MUX2X1 U807 ( .B(n500), .A(n316), .S(n644), .Y(\fifo_next2<5> ) );
  MUX2X1 U808 ( .B(n499), .A(n317), .S(n644), .Y(\fifo_next2<6> ) );
  MUX2X1 U809 ( .B(n498), .A(n318), .S(n644), .Y(\fifo_next2<7> ) );
  MUX2X1 U810 ( .B(n497), .A(n319), .S(n644), .Y(\fifo_next2<8> ) );
  MUX2X1 U811 ( .B(n496), .A(n320), .S(n644), .Y(\fifo_next2<9> ) );
  MUX2X1 U812 ( .B(n495), .A(n321), .S(n644), .Y(\fifo_next2<10> ) );
  MUX2X1 U813 ( .B(n494), .A(n322), .S(n644), .Y(\fifo_next2<11> ) );
  MUX2X1 U814 ( .B(n493), .A(n323), .S(n644), .Y(\fifo_next2<12> ) );
  MUX2X1 U815 ( .B(n492), .A(n324), .S(n643), .Y(\fifo_next2<13> ) );
  MUX2X1 U816 ( .B(n491), .A(n325), .S(n643), .Y(\fifo_next2<14> ) );
  MUX2X1 U817 ( .B(n490), .A(n326), .S(n643), .Y(\fifo_next2<15> ) );
  MUX2X1 U818 ( .B(n489), .A(n327), .S(n643), .Y(\fifo_next2<16> ) );
  MUX2X1 U819 ( .B(n488), .A(n328), .S(n643), .Y(\fifo_next2<17> ) );
  MUX2X1 U820 ( .B(n487), .A(n329), .S(n643), .Y(\fifo_next2<18> ) );
  MUX2X1 U821 ( .B(n486), .A(n330), .S(n643), .Y(\fifo_next2<19> ) );
  MUX2X1 U822 ( .B(n485), .A(n331), .S(n643), .Y(\fifo_next2<20> ) );
  MUX2X1 U823 ( .B(n484), .A(n332), .S(n643), .Y(\fifo_next2<21> ) );
  MUX2X1 U824 ( .B(n483), .A(n333), .S(n643), .Y(\fifo_next2<22> ) );
  MUX2X1 U825 ( .B(n482), .A(n334), .S(n643), .Y(\fifo_next2<23> ) );
  MUX2X1 U826 ( .B(n481), .A(n335), .S(n643), .Y(\fifo_next2<24> ) );
  MUX2X1 U827 ( .B(n480), .A(n336), .S(n644), .Y(\fifo_next2<25> ) );
  MUX2X1 U828 ( .B(n479), .A(n337), .S(n643), .Y(\fifo_next2<26> ) );
  MUX2X1 U829 ( .B(n478), .A(n338), .S(n644), .Y(\fifo_next2<27> ) );
  MUX2X1 U830 ( .B(n477), .A(n339), .S(n643), .Y(\fifo_next2<28> ) );
  MUX2X1 U831 ( .B(n476), .A(n340), .S(n644), .Y(\fifo_next2<29> ) );
  MUX2X1 U832 ( .B(n475), .A(n341), .S(n643), .Y(\fifo_next2<30> ) );
  MUX2X1 U833 ( .B(n474), .A(n342), .S(n644), .Y(\fifo_next2<31> ) );
  MUX2X1 U834 ( .B(n473), .A(n343), .S(n643), .Y(\fifo_next2<32> ) );
  MUX2X1 U835 ( .B(n472), .A(n344), .S(n644), .Y(\fifo_next2<33> ) );
  MUX2X1 U836 ( .B(n471), .A(n345), .S(n643), .Y(\fifo_next2<34> ) );
  MUX2X1 U837 ( .B(n470), .A(n346), .S(n644), .Y(\fifo_next2<35> ) );
  MUX2X1 U838 ( .B(n469), .A(n347), .S(n643), .Y(\fifo_next2<36> ) );
  MUX2X1 U839 ( .B(n468), .A(n348), .S(n642), .Y(\fifo_next2<37> ) );
  MUX2X1 U840 ( .B(n467), .A(n349), .S(n643), .Y(\fifo_next2<38> ) );
  MUX2X1 U841 ( .B(n466), .A(n350), .S(n644), .Y(\fifo_next2<39> ) );
  MUX2X1 U842 ( .B(n465), .A(n351), .S(n642), .Y(\fifo_next2<40> ) );
  MUX2X1 U843 ( .B(n464), .A(n352), .S(n643), .Y(\fifo_next2<41> ) );
  MUX2X1 U844 ( .B(n463), .A(n353), .S(n644), .Y(\fifo_next2<42> ) );
  MUX2X1 U845 ( .B(n462), .A(n354), .S(n642), .Y(\fifo_next2<43> ) );
  MUX2X1 U846 ( .B(n461), .A(n355), .S(n642), .Y(\fifo_next2<44> ) );
  MUX2X1 U847 ( .B(n460), .A(n356), .S(n642), .Y(\fifo_next2<45> ) );
  MUX2X1 U848 ( .B(n459), .A(n357), .S(n642), .Y(\fifo_next2<46> ) );
  MUX2X1 U849 ( .B(n458), .A(n358), .S(n642), .Y(\fifo_next2<47> ) );
  MUX2X1 U850 ( .B(n457), .A(n359), .S(n642), .Y(\fifo_next2<48> ) );
  MUX2X1 U851 ( .B(n456), .A(n360), .S(n642), .Y(\fifo_next2<49> ) );
  MUX2X1 U852 ( .B(n455), .A(n361), .S(n642), .Y(\fifo_next2<50> ) );
  MUX2X1 U853 ( .B(n454), .A(n362), .S(n642), .Y(\fifo_next2<51> ) );
  MUX2X1 U854 ( .B(n453), .A(n363), .S(n642), .Y(\fifo_next2<52> ) );
  MUX2X1 U855 ( .B(n452), .A(n364), .S(n642), .Y(\fifo_next2<53> ) );
  MUX2X1 U856 ( .B(n451), .A(n365), .S(n642), .Y(\fifo_next2<54> ) );
  MUX2X1 U857 ( .B(n450), .A(n366), .S(n642), .Y(\fifo_next2<55> ) );
  MUX2X1 U858 ( .B(n449), .A(n367), .S(n642), .Y(\fifo_next2<56> ) );
  MUX2X1 U859 ( .B(n448), .A(n368), .S(n642), .Y(\fifo_next2<57> ) );
  MUX2X1 U860 ( .B(n447), .A(n369), .S(n642), .Y(\fifo_next2<58> ) );
  MUX2X1 U861 ( .B(n446), .A(n370), .S(n642), .Y(\fifo_next2<59> ) );
  MUX2X1 U862 ( .B(n445), .A(n371), .S(n642), .Y(\fifo_next2<60> ) );
  MUX2X1 U863 ( .B(n444), .A(n372), .S(n644), .Y(\fifo_next2<61> ) );
  MUX2X1 U864 ( .B(n443), .A(n373), .S(n642), .Y(\fifo_next2<62> ) );
  MUX2X1 U865 ( .B(n442), .A(n374), .S(n642), .Y(\fifo_next2<63> ) );
  MUX2X1 U866 ( .B(n569), .A(n311), .S(n296), .Y(\fifo_next1<0> ) );
  MUX2X1 U867 ( .B(n568), .A(n312), .S(n638), .Y(\fifo_next1<1> ) );
  MUX2X1 U868 ( .B(n567), .A(n313), .S(n638), .Y(\fifo_next1<2> ) );
  MUX2X1 U869 ( .B(n566), .A(n314), .S(n638), .Y(\fifo_next1<3> ) );
  MUX2X1 U870 ( .B(n565), .A(n315), .S(n638), .Y(\fifo_next1<4> ) );
  MUX2X1 U871 ( .B(n564), .A(n316), .S(n638), .Y(\fifo_next1<5> ) );
  MUX2X1 U872 ( .B(n563), .A(n317), .S(n638), .Y(\fifo_next1<6> ) );
  MUX2X1 U873 ( .B(n562), .A(n318), .S(n638), .Y(\fifo_next1<7> ) );
  MUX2X1 U874 ( .B(n561), .A(n319), .S(n638), .Y(\fifo_next1<8> ) );
  MUX2X1 U875 ( .B(n560), .A(n320), .S(n638), .Y(\fifo_next1<9> ) );
  MUX2X1 U876 ( .B(n559), .A(n321), .S(n638), .Y(\fifo_next1<10> ) );
  MUX2X1 U877 ( .B(n558), .A(n322), .S(n638), .Y(\fifo_next1<11> ) );
  MUX2X1 U878 ( .B(n557), .A(n323), .S(n638), .Y(\fifo_next1<12> ) );
  MUX2X1 U879 ( .B(n556), .A(n324), .S(n637), .Y(\fifo_next1<13> ) );
  MUX2X1 U880 ( .B(n555), .A(n325), .S(n637), .Y(\fifo_next1<14> ) );
  MUX2X1 U881 ( .B(n554), .A(n326), .S(n637), .Y(\fifo_next1<15> ) );
  MUX2X1 U882 ( .B(n553), .A(n327), .S(n637), .Y(\fifo_next1<16> ) );
  MUX2X1 U883 ( .B(n552), .A(n328), .S(n637), .Y(\fifo_next1<17> ) );
  MUX2X1 U884 ( .B(n551), .A(n329), .S(n637), .Y(\fifo_next1<18> ) );
  MUX2X1 U885 ( .B(n550), .A(n330), .S(n637), .Y(\fifo_next1<19> ) );
  MUX2X1 U886 ( .B(n549), .A(n331), .S(n637), .Y(\fifo_next1<20> ) );
  MUX2X1 U887 ( .B(n548), .A(n332), .S(n637), .Y(\fifo_next1<21> ) );
  MUX2X1 U888 ( .B(n547), .A(n333), .S(n637), .Y(\fifo_next1<22> ) );
  MUX2X1 U889 ( .B(n546), .A(n334), .S(n637), .Y(\fifo_next1<23> ) );
  MUX2X1 U890 ( .B(n545), .A(n335), .S(n637), .Y(\fifo_next1<24> ) );
  MUX2X1 U891 ( .B(n544), .A(n336), .S(n637), .Y(\fifo_next1<25> ) );
  MUX2X1 U892 ( .B(n543), .A(n337), .S(n638), .Y(\fifo_next1<26> ) );
  MUX2X1 U893 ( .B(n542), .A(n338), .S(n637), .Y(\fifo_next1<27> ) );
  MUX2X1 U894 ( .B(n541), .A(n339), .S(n638), .Y(\fifo_next1<28> ) );
  MUX2X1 U895 ( .B(n540), .A(n340), .S(n637), .Y(\fifo_next1<29> ) );
  MUX2X1 U896 ( .B(n539), .A(n341), .S(n638), .Y(\fifo_next1<30> ) );
  MUX2X1 U897 ( .B(n538), .A(n342), .S(n637), .Y(\fifo_next1<31> ) );
  MUX2X1 U898 ( .B(n537), .A(n343), .S(n638), .Y(\fifo_next1<32> ) );
  MUX2X1 U899 ( .B(n536), .A(n344), .S(n637), .Y(\fifo_next1<33> ) );
  MUX2X1 U900 ( .B(n535), .A(n345), .S(n638), .Y(\fifo_next1<34> ) );
  MUX2X1 U901 ( .B(n534), .A(n346), .S(n637), .Y(\fifo_next1<35> ) );
  MUX2X1 U902 ( .B(n533), .A(n347), .S(n638), .Y(\fifo_next1<36> ) );
  MUX2X1 U903 ( .B(n532), .A(n348), .S(n636), .Y(\fifo_next1<37> ) );
  MUX2X1 U904 ( .B(n531), .A(n349), .S(n636), .Y(\fifo_next1<38> ) );
  MUX2X1 U905 ( .B(n530), .A(n350), .S(n636), .Y(\fifo_next1<39> ) );
  MUX2X1 U906 ( .B(n529), .A(n351), .S(n636), .Y(\fifo_next1<40> ) );
  MUX2X1 U907 ( .B(n528), .A(n352), .S(n636), .Y(\fifo_next1<41> ) );
  MUX2X1 U908 ( .B(n527), .A(n353), .S(n636), .Y(\fifo_next1<42> ) );
  MUX2X1 U909 ( .B(n526), .A(n354), .S(n636), .Y(\fifo_next1<43> ) );
  MUX2X1 U910 ( .B(n525), .A(n355), .S(n636), .Y(\fifo_next1<44> ) );
  MUX2X1 U911 ( .B(n524), .A(n356), .S(n636), .Y(\fifo_next1<45> ) );
  MUX2X1 U912 ( .B(n523), .A(n357), .S(n636), .Y(\fifo_next1<46> ) );
  MUX2X1 U913 ( .B(n522), .A(n358), .S(n636), .Y(\fifo_next1<47> ) );
  MUX2X1 U914 ( .B(n521), .A(n359), .S(n636), .Y(\fifo_next1<48> ) );
  MUX2X1 U915 ( .B(n520), .A(n360), .S(n637), .Y(\fifo_next1<49> ) );
  MUX2X1 U916 ( .B(n519), .A(n361), .S(n636), .Y(\fifo_next1<50> ) );
  MUX2X1 U917 ( .B(n518), .A(n362), .S(n638), .Y(\fifo_next1<51> ) );
  MUX2X1 U918 ( .B(n517), .A(n363), .S(n637), .Y(\fifo_next1<52> ) );
  MUX2X1 U919 ( .B(n516), .A(n364), .S(n636), .Y(\fifo_next1<53> ) );
  MUX2X1 U920 ( .B(n515), .A(n365), .S(n638), .Y(\fifo_next1<54> ) );
  MUX2X1 U921 ( .B(n514), .A(n366), .S(n637), .Y(\fifo_next1<55> ) );
  MUX2X1 U922 ( .B(n513), .A(n367), .S(n636), .Y(\fifo_next1<56> ) );
  MUX2X1 U923 ( .B(n512), .A(n368), .S(n636), .Y(\fifo_next1<57> ) );
  MUX2X1 U924 ( .B(n511), .A(n369), .S(n636), .Y(\fifo_next1<58> ) );
  MUX2X1 U925 ( .B(n510), .A(n370), .S(n636), .Y(\fifo_next1<59> ) );
  MUX2X1 U926 ( .B(n509), .A(n371), .S(n636), .Y(\fifo_next1<60> ) );
  MUX2X1 U927 ( .B(n508), .A(n372), .S(n636), .Y(\fifo_next1<61> ) );
  MUX2X1 U928 ( .B(n507), .A(n373), .S(n636), .Y(\fifo_next1<62> ) );
  MUX2X1 U929 ( .B(n506), .A(n374), .S(n636), .Y(\fifo_next1<63> ) );
  MUX2X1 U930 ( .B(n375), .A(n311), .S(n298), .Y(\fifo_next0<0> ) );
  MUX2X1 U931 ( .B(n632), .A(n312), .S(n641), .Y(\fifo_next0<1> ) );
  MUX2X1 U932 ( .B(n631), .A(n313), .S(n641), .Y(\fifo_next0<2> ) );
  MUX2X1 U933 ( .B(n630), .A(n314), .S(n641), .Y(\fifo_next0<3> ) );
  MUX2X1 U934 ( .B(n629), .A(n315), .S(n641), .Y(\fifo_next0<4> ) );
  MUX2X1 U935 ( .B(n628), .A(n316), .S(n641), .Y(\fifo_next0<5> ) );
  MUX2X1 U936 ( .B(n627), .A(n317), .S(n641), .Y(\fifo_next0<6> ) );
  MUX2X1 U937 ( .B(n626), .A(n318), .S(n641), .Y(\fifo_next0<7> ) );
  MUX2X1 U938 ( .B(n625), .A(n319), .S(n641), .Y(\fifo_next0<8> ) );
  MUX2X1 U939 ( .B(n624), .A(n320), .S(n641), .Y(\fifo_next0<9> ) );
  MUX2X1 U940 ( .B(n623), .A(n321), .S(n641), .Y(\fifo_next0<10> ) );
  MUX2X1 U941 ( .B(n622), .A(n322), .S(n641), .Y(\fifo_next0<11> ) );
  MUX2X1 U942 ( .B(n621), .A(n323), .S(n641), .Y(\fifo_next0<12> ) );
  MUX2X1 U943 ( .B(n620), .A(n324), .S(n640), .Y(\fifo_next0<13> ) );
  MUX2X1 U944 ( .B(n619), .A(n325), .S(n640), .Y(\fifo_next0<14> ) );
  MUX2X1 U945 ( .B(n618), .A(n326), .S(n640), .Y(\fifo_next0<15> ) );
  MUX2X1 U946 ( .B(n617), .A(n327), .S(n640), .Y(\fifo_next0<16> ) );
  MUX2X1 U947 ( .B(n616), .A(n328), .S(n640), .Y(\fifo_next0<17> ) );
  MUX2X1 U948 ( .B(n615), .A(n329), .S(n640), .Y(\fifo_next0<18> ) );
  MUX2X1 U949 ( .B(n614), .A(n330), .S(n640), .Y(\fifo_next0<19> ) );
  MUX2X1 U950 ( .B(n613), .A(n331), .S(n640), .Y(\fifo_next0<20> ) );
  MUX2X1 U951 ( .B(n612), .A(n332), .S(n640), .Y(\fifo_next0<21> ) );
  MUX2X1 U952 ( .B(n611), .A(n333), .S(n640), .Y(\fifo_next0<22> ) );
  MUX2X1 U953 ( .B(n610), .A(n334), .S(n640), .Y(\fifo_next0<23> ) );
  MUX2X1 U954 ( .B(n609), .A(n335), .S(n640), .Y(\fifo_next0<24> ) );
  MUX2X1 U955 ( .B(n608), .A(n336), .S(n640), .Y(\fifo_next0<25> ) );
  MUX2X1 U956 ( .B(n607), .A(n337), .S(n641), .Y(\fifo_next0<26> ) );
  MUX2X1 U957 ( .B(n606), .A(n338), .S(n640), .Y(\fifo_next0<27> ) );
  MUX2X1 U958 ( .B(n605), .A(n339), .S(n641), .Y(\fifo_next0<28> ) );
  MUX2X1 U959 ( .B(n604), .A(n340), .S(n640), .Y(\fifo_next0<29> ) );
  MUX2X1 U960 ( .B(n603), .A(n341), .S(n641), .Y(\fifo_next0<30> ) );
  MUX2X1 U961 ( .B(n602), .A(n342), .S(n640), .Y(\fifo_next0<31> ) );
  MUX2X1 U962 ( .B(n601), .A(n343), .S(n641), .Y(\fifo_next0<32> ) );
  MUX2X1 U963 ( .B(n600), .A(n344), .S(n640), .Y(\fifo_next0<33> ) );
  MUX2X1 U964 ( .B(n599), .A(n345), .S(n641), .Y(\fifo_next0<34> ) );
  MUX2X1 U965 ( .B(n598), .A(n346), .S(n640), .Y(\fifo_next0<35> ) );
  MUX2X1 U966 ( .B(n597), .A(n347), .S(n641), .Y(\fifo_next0<36> ) );
  MUX2X1 U967 ( .B(n596), .A(n348), .S(n639), .Y(\fifo_next0<37> ) );
  MUX2X1 U968 ( .B(n595), .A(n349), .S(n639), .Y(\fifo_next0<38> ) );
  MUX2X1 U969 ( .B(n594), .A(n350), .S(n639), .Y(\fifo_next0<39> ) );
  MUX2X1 U970 ( .B(n593), .A(n351), .S(n639), .Y(\fifo_next0<40> ) );
  MUX2X1 U971 ( .B(n592), .A(n352), .S(n639), .Y(\fifo_next0<41> ) );
  MUX2X1 U972 ( .B(n591), .A(n353), .S(n639), .Y(\fifo_next0<42> ) );
  MUX2X1 U973 ( .B(n590), .A(n354), .S(n639), .Y(\fifo_next0<43> ) );
  MUX2X1 U974 ( .B(n589), .A(n355), .S(n639), .Y(\fifo_next0<44> ) );
  MUX2X1 U975 ( .B(n588), .A(n356), .S(n639), .Y(\fifo_next0<45> ) );
  MUX2X1 U976 ( .B(n587), .A(n357), .S(n639), .Y(\fifo_next0<46> ) );
  MUX2X1 U977 ( .B(n586), .A(n358), .S(n639), .Y(\fifo_next0<47> ) );
  MUX2X1 U978 ( .B(n585), .A(n359), .S(n639), .Y(\fifo_next0<48> ) );
  MUX2X1 U979 ( .B(n584), .A(n360), .S(n640), .Y(\fifo_next0<49> ) );
  MUX2X1 U980 ( .B(n583), .A(n361), .S(n639), .Y(\fifo_next0<50> ) );
  MUX2X1 U981 ( .B(n582), .A(n362), .S(n641), .Y(\fifo_next0<51> ) );
  MUX2X1 U982 ( .B(n581), .A(n363), .S(n640), .Y(\fifo_next0<52> ) );
  MUX2X1 U983 ( .B(n580), .A(n364), .S(n639), .Y(\fifo_next0<53> ) );
  MUX2X1 U984 ( .B(n579), .A(n365), .S(n641), .Y(\fifo_next0<54> ) );
  MUX2X1 U985 ( .B(n578), .A(n366), .S(n640), .Y(\fifo_next0<55> ) );
  MUX2X1 U986 ( .B(n577), .A(n367), .S(n639), .Y(\fifo_next0<56> ) );
  MUX2X1 U987 ( .B(n576), .A(n368), .S(n639), .Y(\fifo_next0<57> ) );
  MUX2X1 U988 ( .B(n575), .A(n369), .S(n639), .Y(\fifo_next0<58> ) );
  MUX2X1 U989 ( .B(n574), .A(n370), .S(n639), .Y(\fifo_next0<59> ) );
  MUX2X1 U990 ( .B(n573), .A(n371), .S(n639), .Y(\fifo_next0<60> ) );
  MUX2X1 U991 ( .B(n572), .A(n372), .S(n639), .Y(\fifo_next0<61> ) );
  MUX2X1 U992 ( .B(n571), .A(n373), .S(n639), .Y(\fifo_next0<62> ) );
  MUX2X1 U993 ( .B(n570), .A(n374), .S(n639), .Y(\fifo_next0<63> ) );
  NAND3X1 U994 ( .A(\writestate<1> ), .B(n306), .C(\writestate<0> ), .Y(n307)
         );
  NAND3X1 U995 ( .A(n306), .B(n377), .C(\writestate<1> ), .Y(n308) );
  NAND3X1 U996 ( .A(n306), .B(n376), .C(\writestate<0> ), .Y(n309) );
  NAND3X1 U997 ( .A(n376), .B(n377), .C(n306), .Y(n310) );
endmodule

