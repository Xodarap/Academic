library verilog;
use verilog.vl_types.all;
entity tb_rf is
end tb_rf;
