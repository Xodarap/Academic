library verilog;
use verilog.vl_types.all;
entity mem_system_perfbench is
end mem_system_perfbench;
