library verilog;
use verilog.vl_types.all;
entity tb_add2 is
end tb_add2;
