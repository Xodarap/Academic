library verilog;
use verilog.vl_types.all;
entity tb_adder16 is
end tb_adder16;
