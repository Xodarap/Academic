library verilog;
use verilog.vl_types.all;
entity proc_hier_bench is
end proc_hier_bench;
