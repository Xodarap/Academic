library verilog;
use verilog.vl_types.all;
entity tb_decode is
end tb_decode;
