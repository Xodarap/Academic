library verilog;
use verilog.vl_types.all;
entity rf_bench is
end rf_bench;
