library verilog;
use verilog.vl_types.all;
entity mem_interface_tb is
end mem_interface_tb;
